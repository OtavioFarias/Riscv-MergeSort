`timescale 1ns/1ps

module tb_top;

  reg clk;
  reg reset;

  // Instância do módulo top
  Top uut (
    .realClock(clk),
    .reset(reset)
  );

  initial begin
    // Geração do VCD
    $dumpfile("projeto/build/dump.vcd");
    $dumpvars(0, tb_top);

    // Inicialização dos sinais
    clk = 0;
    reset = 1;

    // Aguarda 20ns com reset ativo
    #20;
    reset = 0;

    // Roda a simulação por mais 200ns
    //#16499280;
    #20_000_000;
    //#62_914_560;

    // Finaliza a simulação
    $finish;
  end

  // Geração de clock (10ns de período: 5ns alto, 5ns baixo)
  always #5 clk = ~clk;

endmodule

module RAM(

    input [31:0] address,
    input [31:0] value,
    output [31:0] data,
    input write,
    input clock,
    output stallSignal,
	input read,
	input reset
);

reg [7:0] memory[0:32000];

initial begin

    $readmemb("projeto/dadosUnificados1024.txt", memory);

end

reg [1:0] stall;

assign stallSignal = (stall == 2'b11) ? 1'b1 : 1'b0;
//assign stallSignal = 1'b0;



assign data = {memory[address], memory[address+1], memory[address+2], memory[address+3]};

always @(posedge clock, posedge reset) begin

	if(reset) begin

		stall <= 2'b0;

	end
	else begin

		stall <= stall + 1;

		if(write) begin

		    memory[address] = value[31:24];
		    memory[address + 1] = value[23:16];
		    memory[address + 2] = value[15:8];
		    memory[address + 3] = value[7:0];

		end
	end
end

wire [31:0] memory0 = {memory[0], memory[1], memory[2], memory[3]};
wire [31:0] memory4 = {memory[4], memory[5], memory[6], memory[7]};
wire [31:0] memory8 = {memory[8], memory[9], memory[10], memory[11]};
wire [31:0] memory12 = {memory[12], memory[13], memory[14], memory[15]};
wire [31:0] memory16 = {memory[16], memory[17], memory[18], memory[19]};
wire [31:0] memory20 = {memory[20], memory[21], memory[22], memory[23]};
wire [31:0] memory24 = {memory[24], memory[25], memory[26], memory[27]};
wire [31:0] memory28 = {memory[28], memory[29], memory[30], memory[31]};
wire [31:0] memory32 = {memory[32], memory[33], memory[34], memory[35]};
wire [31:0] memory36 = {memory[36], memory[37], memory[38], memory[39]};
wire [31:0] memory40 = {memory[40], memory[41], memory[42], memory[43]};
wire [31:0] memory44 = {memory[44], memory[45], memory[46], memory[47]};
wire [31:0] memory48 = {memory[48], memory[49], memory[50], memory[51]};
wire [31:0] memory52 = {memory[52], memory[53], memory[54], memory[55]};
wire [31:0] memory56 = {memory[56], memory[57], memory[58], memory[59]};
wire [31:0] memory60 = {memory[60], memory[61], memory[62], memory[63]};
wire [31:0] memory64 = {memory[64], memory[65], memory[66], memory[67]};
wire [31:0] memory68 = {memory[68], memory[69], memory[70], memory[71]};
wire [31:0] memory72 = {memory[72], memory[73], memory[74], memory[75]};
wire [31:0] memory76 = {memory[76], memory[77], memory[78], memory[79]};
wire [31:0] memory80 = {memory[80], memory[81], memory[82], memory[83]};
wire [31:0] memory84 = {memory[84], memory[85], memory[86], memory[87]};
wire [31:0] memory88 = {memory[88], memory[89], memory[90], memory[91]};
wire [31:0] memory92 = {memory[92], memory[93], memory[94], memory[95]};
wire [31:0] memory96 = {memory[96], memory[97], memory[98], memory[99]};
wire [31:0] memory100 = {memory[100], memory[101], memory[102], memory[103]};
wire [31:0] memory104 = {memory[104], memory[105], memory[106], memory[107]};
wire [31:0] memory108 = {memory[108], memory[109], memory[110], memory[111]};
wire [31:0] memory112 = {memory[112], memory[113], memory[114], memory[115]};
wire [31:0] memory116 = {memory[116], memory[117], memory[118], memory[119]};
wire [31:0] memory120 = {memory[120], memory[121], memory[122], memory[123]};
wire [31:0] memory124 = {memory[124], memory[125], memory[126], memory[127]};
wire [31:0] memory128 = {memory[128], memory[129], memory[130], memory[131]};
wire [31:0] memory132 = {memory[132], memory[133], memory[134], memory[135]};
wire [31:0] memory136 = {memory[136], memory[137], memory[138], memory[139]};
wire [31:0] memory140 = {memory[140], memory[141], memory[142], memory[143]};
wire [31:0] memory144 = {memory[144], memory[145], memory[146], memory[147]};
wire [31:0] memory148 = {memory[148], memory[149], memory[150], memory[151]};
wire [31:0] memory152 = {memory[152], memory[153], memory[154], memory[155]};
wire [31:0] memory156 = {memory[156], memory[157], memory[158], memory[159]};
wire [31:0] memory160 = {memory[160], memory[161], memory[162], memory[163]};
wire [31:0] memory164 = {memory[164], memory[165], memory[166], memory[167]};
wire [31:0] memory168 = {memory[168], memory[169], memory[170], memory[171]};
wire [31:0] memory172 = {memory[172], memory[173], memory[174], memory[175]};
wire [31:0] memory176 = {memory[176], memory[177], memory[178], memory[179]};
wire [31:0] memory180 = {memory[180], memory[181], memory[182], memory[183]};
wire [31:0] memory184 = {memory[184], memory[185], memory[186], memory[187]};
wire [31:0] memory188 = {memory[188], memory[189], memory[190], memory[191]};
wire [31:0] memory192 = {memory[192], memory[193], memory[194], memory[195]};
wire [31:0] memory196 = {memory[196], memory[197], memory[198], memory[199]};
wire [31:0] memory200 = {memory[200], memory[201], memory[202], memory[203]};
wire [31:0] memory204 = {memory[204], memory[205], memory[206], memory[207]};
wire [31:0] memory208 = {memory[208], memory[209], memory[210], memory[211]};
wire [31:0] memory212 = {memory[212], memory[213], memory[214], memory[215]};
wire [31:0] memory216 = {memory[216], memory[217], memory[218], memory[219]};
wire [31:0] memory220 = {memory[220], memory[221], memory[222], memory[223]};
wire [31:0] memory224 = {memory[224], memory[225], memory[226], memory[227]};
wire [31:0] memory228 = {memory[228], memory[229], memory[230], memory[231]};
wire [31:0] memory232 = {memory[232], memory[233], memory[234], memory[235]};
wire [31:0] memory236 = {memory[236], memory[237], memory[238], memory[239]};
wire [31:0] memory240 = {memory[240], memory[241], memory[242], memory[243]};
wire [31:0] memory244 = {memory[244], memory[245], memory[246], memory[247]};
wire [31:0] memory248 = {memory[248], memory[249], memory[250], memory[251]};
wire [31:0] memory252 = {memory[252], memory[253], memory[254], memory[255]};
wire [31:0] memory256 = {memory[256], memory[257], memory[258], memory[259]};
wire [31:0] memory260 = {memory[260], memory[261], memory[262], memory[263]};
wire [31:0] memory264 = {memory[264], memory[265], memory[266], memory[267]};
wire [31:0] memory268 = {memory[268], memory[269], memory[270], memory[271]};
wire [31:0] memory272 = {memory[272], memory[273], memory[274], memory[275]};
wire [31:0] memory276 = {memory[276], memory[277], memory[278], memory[279]};
wire [31:0] memory280 = {memory[280], memory[281], memory[282], memory[283]};
wire [31:0] memory284 = {memory[284], memory[285], memory[286], memory[287]};
wire [31:0] memory288 = {memory[288], memory[289], memory[290], memory[291]};
wire [31:0] memory292 = {memory[292], memory[293], memory[294], memory[295]};
wire [31:0] memory296 = {memory[296], memory[297], memory[298], memory[299]};
wire [31:0] memory300 = {memory[300], memory[301], memory[302], memory[303]};
wire [31:0] memory304 = {memory[304], memory[305], memory[306], memory[307]};
wire [31:0] memory308 = {memory[308], memory[309], memory[310], memory[311]};
wire [31:0] memory312 = {memory[312], memory[313], memory[314], memory[315]};
wire [31:0] memory316 = {memory[316], memory[317], memory[318], memory[319]};
wire [31:0] memory320 = {memory[320], memory[321], memory[322], memory[323]};
wire [31:0] memory324 = {memory[324], memory[325], memory[326], memory[327]};
wire [31:0] memory328 = {memory[328], memory[329], memory[330], memory[331]};
wire [31:0] memory332 = {memory[332], memory[333], memory[334], memory[335]};
wire [31:0] memory336 = {memory[336], memory[337], memory[338], memory[339]};
wire [31:0] memory340 = {memory[340], memory[341], memory[342], memory[343]};
wire [31:0] memory344 = {memory[344], memory[345], memory[346], memory[347]};
wire [31:0] memory348 = {memory[348], memory[349], memory[350], memory[351]};
wire [31:0] memory352 = {memory[352], memory[353], memory[354], memory[355]};
wire [31:0] memory356 = {memory[356], memory[357], memory[358], memory[359]};
wire [31:0] memory360 = {memory[360], memory[361], memory[362], memory[363]};
wire [31:0] memory364 = {memory[364], memory[365], memory[366], memory[367]};
wire [31:0] memory368 = {memory[368], memory[369], memory[370], memory[371]};
wire [31:0] memory372 = {memory[372], memory[373], memory[374], memory[375]};
wire [31:0] memory376 = {memory[376], memory[377], memory[378], memory[379]};
wire [31:0] memory380 = {memory[380], memory[381], memory[382], memory[383]};
wire [31:0] memory384 = {memory[384], memory[385], memory[386], memory[387]};
wire [31:0] memory388 = {memory[388], memory[389], memory[390], memory[391]};
wire [31:0] memory392 = {memory[392], memory[393], memory[394], memory[395]};
wire [31:0] memory396 = {memory[396], memory[397], memory[398], memory[399]};
wire [31:0] memory400 = {memory[400], memory[401], memory[402], memory[403]};
wire [31:0] memory404 = {memory[404], memory[405], memory[406], memory[407]};
wire [31:0] memory408 = {memory[408], memory[409], memory[410], memory[411]};
wire [31:0] memory412 = {memory[412], memory[413], memory[414], memory[415]};
wire [31:0] memory416 = {memory[416], memory[417], memory[418], memory[419]};
wire [31:0] memory420 = {memory[420], memory[421], memory[422], memory[423]};
wire [31:0] memory424 = {memory[424], memory[425], memory[426], memory[427]};
wire [31:0] memory428 = {memory[428], memory[429], memory[430], memory[431]};
wire [31:0] memory432 = {memory[432], memory[433], memory[434], memory[435]};
wire [31:0] memory436 = {memory[436], memory[437], memory[438], memory[439]};
wire [31:0] memory440 = {memory[440], memory[441], memory[442], memory[443]};
wire [31:0] memory444 = {memory[444], memory[445], memory[446], memory[447]};
wire [31:0] memory448 = {memory[448], memory[449], memory[450], memory[451]};
wire [31:0] memory452 = {memory[452], memory[453], memory[454], memory[455]};
wire [31:0] memory456 = {memory[456], memory[457], memory[458], memory[459]};
wire [31:0] memory460 = {memory[460], memory[461], memory[462], memory[463]};
wire [31:0] memory464 = {memory[464], memory[465], memory[466], memory[467]};
wire [31:0] memory468 = {memory[468], memory[469], memory[470], memory[471]};
wire [31:0] memory472 = {memory[472], memory[473], memory[474], memory[475]};
wire [31:0] memory476 = {memory[476], memory[477], memory[478], memory[479]};
wire [31:0] memory480 = {memory[480], memory[481], memory[482], memory[483]};
wire [31:0] memory484 = {memory[484], memory[485], memory[486], memory[487]};
wire [31:0] memory488 = {memory[488], memory[489], memory[490], memory[491]};
wire [31:0] memory492 = {memory[492], memory[493], memory[494], memory[495]};
wire [31:0] memory496 = {memory[496], memory[497], memory[498], memory[499]};
wire [31:0] memory500 = {memory[500], memory[501], memory[502], memory[503]};
wire [31:0] memory504 = {memory[504], memory[505], memory[506], memory[507]};
wire [31:0] memory508 = {memory[508], memory[509], memory[510], memory[511]};
wire [31:0] memory512 = {memory[512], memory[513], memory[514], memory[515]};
wire [31:0] memory516 = {memory[516], memory[517], memory[518], memory[519]};
wire [31:0] memory520 = {memory[520], memory[521], memory[522], memory[523]};
wire [31:0] memory524 = {memory[524], memory[525], memory[526], memory[527]};
wire [31:0] memory528 = {memory[528], memory[529], memory[530], memory[531]};
wire [31:0] memory532 = {memory[532], memory[533], memory[534], memory[535]};
wire [31:0] memory536 = {memory[536], memory[537], memory[538], memory[539]};
wire [31:0] memory540 = {memory[540], memory[541], memory[542], memory[543]};
wire [31:0] memory544 = {memory[544], memory[545], memory[546], memory[547]};
wire [31:0] memory548 = {memory[548], memory[549], memory[550], memory[551]};
wire [31:0] memory552 = {memory[552], memory[553], memory[554], memory[555]};
wire [31:0] memory556 = {memory[556], memory[557], memory[558], memory[559]};
wire [31:0] memory560 = {memory[560], memory[561], memory[562], memory[563]};
wire [31:0] memory564 = {memory[564], memory[565], memory[566], memory[567]};
wire [31:0] memory568 = {memory[568], memory[569], memory[570], memory[571]};
wire [31:0] memory572 = {memory[572], memory[573], memory[574], memory[575]};
wire [31:0] memory576 = {memory[576], memory[577], memory[578], memory[579]};
wire [31:0] memory580 = {memory[580], memory[581], memory[582], memory[583]};
wire [31:0] memory584 = {memory[584], memory[585], memory[586], memory[587]};
wire [31:0] memory588 = {memory[588], memory[589], memory[590], memory[591]};
wire [31:0] memory592 = {memory[592], memory[593], memory[594], memory[595]};
wire [31:0] memory596 = {memory[596], memory[597], memory[598], memory[599]};
wire [31:0] memory600 = {memory[600], memory[601], memory[602], memory[603]};
wire [31:0] memory604 = {memory[604], memory[605], memory[606], memory[607]};
wire [31:0] memory608 = {memory[608], memory[609], memory[610], memory[611]};
wire [31:0] memory612 = {memory[612], memory[613], memory[614], memory[615]};
wire [31:0] memory616 = {memory[616], memory[617], memory[618], memory[619]};
wire [31:0] memory620 = {memory[620], memory[621], memory[622], memory[623]};
wire [31:0] memory624 = {memory[624], memory[625], memory[626], memory[627]};
wire [31:0] memory628 = {memory[628], memory[629], memory[630], memory[631]};
wire [31:0] memory632 = {memory[632], memory[633], memory[634], memory[635]};
wire [31:0] memory636 = {memory[636], memory[637], memory[638], memory[639]};
wire [31:0] memory640 = {memory[640], memory[641], memory[642], memory[643]};
wire [31:0] memory644 = {memory[644], memory[645], memory[646], memory[647]};
wire [31:0] memory648 = {memory[648], memory[649], memory[650], memory[651]};
wire [31:0] memory652 = {memory[652], memory[653], memory[654], memory[655]};
wire [31:0] memory656 = {memory[656], memory[657], memory[658], memory[659]};
wire [31:0] memory660 = {memory[660], memory[661], memory[662], memory[663]};
wire [31:0] memory664 = {memory[664], memory[665], memory[666], memory[667]};
wire [31:0] memory668 = {memory[668], memory[669], memory[670], memory[671]};
wire [31:0] memory672 = {memory[672], memory[673], memory[674], memory[675]};
wire [31:0] memory676 = {memory[676], memory[677], memory[678], memory[679]};
wire [31:0] memory680 = {memory[680], memory[681], memory[682], memory[683]};
wire [31:0] memory684 = {memory[684], memory[685], memory[686], memory[687]};
wire [31:0] memory688 = {memory[688], memory[689], memory[690], memory[691]};
wire [31:0] memory692 = {memory[692], memory[693], memory[694], memory[695]};
wire [31:0] memory696 = {memory[696], memory[697], memory[698], memory[699]};
wire [31:0] memory700 = {memory[700], memory[701], memory[702], memory[703]};
wire [31:0] memory704 = {memory[704], memory[705], memory[706], memory[707]};
wire [31:0] memory708 = {memory[708], memory[709], memory[710], memory[711]};
wire [31:0] memory712 = {memory[712], memory[713], memory[714], memory[715]};
wire [31:0] memory716 = {memory[716], memory[717], memory[718], memory[719]};
wire [31:0] memory720 = {memory[720], memory[721], memory[722], memory[723]};
wire [31:0] memory724 = {memory[724], memory[725], memory[726], memory[727]};
wire [31:0] memory728 = {memory[728], memory[729], memory[730], memory[731]};
wire [31:0] memory732 = {memory[732], memory[733], memory[734], memory[735]};
wire [31:0] memory736 = {memory[736], memory[737], memory[738], memory[739]};
wire [31:0] memory740 = {memory[740], memory[741], memory[742], memory[743]};
wire [31:0] memory744 = {memory[744], memory[745], memory[746], memory[747]};
wire [31:0] memory748 = {memory[748], memory[749], memory[750], memory[751]};
wire [31:0] memory752 = {memory[752], memory[753], memory[754], memory[755]};
wire [31:0] memory756 = {memory[756], memory[757], memory[758], memory[759]};
wire [31:0] memory760 = {memory[760], memory[761], memory[762], memory[763]};
wire [31:0] memory764 = {memory[764], memory[765], memory[766], memory[767]};
wire [31:0] memory768 = {memory[768], memory[769], memory[770], memory[771]};
wire [31:0] memory772 = {memory[772], memory[773], memory[774], memory[775]};
wire [31:0] memory776 = {memory[776], memory[777], memory[778], memory[779]};
wire [31:0] memory780 = {memory[780], memory[781], memory[782], memory[783]};
wire [31:0] memory784 = {memory[784], memory[785], memory[786], memory[787]};
wire [31:0] memory788 = {memory[788], memory[789], memory[790], memory[791]};
wire [31:0] memory792 = {memory[792], memory[793], memory[794], memory[795]};
wire [31:0] memory796 = {memory[796], memory[797], memory[798], memory[799]};
wire [31:0] memory800 = {memory[800], memory[801], memory[802], memory[803]};
wire [31:0] memory804 = {memory[804], memory[805], memory[806], memory[807]};
wire [31:0] memory808 = {memory[808], memory[809], memory[810], memory[811]};
wire [31:0] memory812 = {memory[812], memory[813], memory[814], memory[815]};
wire [31:0] memory816 = {memory[816], memory[817], memory[818], memory[819]};
wire [31:0] memory820 = {memory[820], memory[821], memory[822], memory[823]};
wire [31:0] memory824 = {memory[824], memory[825], memory[826], memory[827]};
wire [31:0] memory828 = {memory[828], memory[829], memory[830], memory[831]};
wire [31:0] memory832 = {memory[832], memory[833], memory[834], memory[835]};
wire [31:0] memory836 = {memory[836], memory[837], memory[838], memory[839]};
wire [31:0] memory840 = {memory[840], memory[841], memory[842], memory[843]};
wire [31:0] memory844 = {memory[844], memory[845], memory[846], memory[847]};
wire [31:0] memory848 = {memory[848], memory[849], memory[850], memory[851]};
wire [31:0] memory852 = {memory[852], memory[853], memory[854], memory[855]};
wire [31:0] memory856 = {memory[856], memory[857], memory[858], memory[859]};
wire [31:0] memory860 = {memory[860], memory[861], memory[862], memory[863]};
wire [31:0] memory864 = {memory[864], memory[865], memory[866], memory[867]};
wire [31:0] memory868 = {memory[868], memory[869], memory[870], memory[871]};
wire [31:0] memory872 = {memory[872], memory[873], memory[874], memory[875]};
wire [31:0] memory876 = {memory[876], memory[877], memory[878], memory[879]};
wire [31:0] memory880 = {memory[880], memory[881], memory[882], memory[883]};
wire [31:0] memory884 = {memory[884], memory[885], memory[886], memory[887]};
wire [31:0] memory888 = {memory[888], memory[889], memory[890], memory[891]};
wire [31:0] memory892 = {memory[892], memory[893], memory[894], memory[895]};
wire [31:0] memory896 = {memory[896], memory[897], memory[898], memory[899]};
wire [31:0] memory900 = {memory[900], memory[901], memory[902], memory[903]};
wire [31:0] memory904 = {memory[904], memory[905], memory[906], memory[907]};
wire [31:0] memory908 = {memory[908], memory[909], memory[910], memory[911]};
wire [31:0] memory912 = {memory[912], memory[913], memory[914], memory[915]};
wire [31:0] memory916 = {memory[916], memory[917], memory[918], memory[919]};
wire [31:0] memory920 = {memory[920], memory[921], memory[922], memory[923]};
wire [31:0] memory924 = {memory[924], memory[925], memory[926], memory[927]};
wire [31:0] memory928 = {memory[928], memory[929], memory[930], memory[931]};
wire [31:0] memory932 = {memory[932], memory[933], memory[934], memory[935]};
wire [31:0] memory936 = {memory[936], memory[937], memory[938], memory[939]};
wire [31:0] memory940 = {memory[940], memory[941], memory[942], memory[943]};
wire [31:0] memory944 = {memory[944], memory[945], memory[946], memory[947]};
wire [31:0] memory948 = {memory[948], memory[949], memory[950], memory[951]};
wire [31:0] memory952 = {memory[952], memory[953], memory[954], memory[955]};
wire [31:0] memory956 = {memory[956], memory[957], memory[958], memory[959]};
wire [31:0] memory960 = {memory[960], memory[961], memory[962], memory[963]};
wire [31:0] memory964 = {memory[964], memory[965], memory[966], memory[967]};
wire [31:0] memory968 = {memory[968], memory[969], memory[970], memory[971]};
wire [31:0] memory972 = {memory[972], memory[973], memory[974], memory[975]};
wire [31:0] memory976 = {memory[976], memory[977], memory[978], memory[979]};
wire [31:0] memory980 = {memory[980], memory[981], memory[982], memory[983]};
wire [31:0] memory984 = {memory[984], memory[985], memory[986], memory[987]};
wire [31:0] memory988 = {memory[988], memory[989], memory[990], memory[991]};
wire [31:0] memory992 = {memory[992], memory[993], memory[994], memory[995]};
wire [31:0] memory996 = {memory[996], memory[997], memory[998], memory[999]};
wire [31:0] memory1000 = {memory[1000], memory[1001], memory[1002], memory[1003]};
wire [31:0] memory1004 = {memory[1004], memory[1005], memory[1006], memory[1007]};
wire [31:0] memory1008 = {memory[1008], memory[1009], memory[1010], memory[1011]};
wire [31:0] memory1012 = {memory[1012], memory[1013], memory[1014], memory[1015]};
wire [31:0] memory1016 = {memory[1016], memory[1017], memory[1018], memory[1019]};
wire [31:0] memory1020 = {memory[1020], memory[1021], memory[1022], memory[1023]};
wire [31:0] memory1024 = {memory[1024], memory[1025], memory[1026], memory[1027]};
wire [31:0] memory1028 = {memory[1028], memory[1029], memory[1030], memory[1031]};
wire [31:0] memory1032 = {memory[1032], memory[1033], memory[1034], memory[1035]};
wire [31:0] memory1036 = {memory[1036], memory[1037], memory[1038], memory[1039]};
wire [31:0] memory1040 = {memory[1040], memory[1041], memory[1042], memory[1043]};
wire [31:0] memory1044 = {memory[1044], memory[1045], memory[1046], memory[1047]};
wire [31:0] memory1048 = {memory[1048], memory[1049], memory[1050], memory[1051]};
wire [31:0] memory1052 = {memory[1052], memory[1053], memory[1054], memory[1055]};
wire [31:0] memory1056 = {memory[1056], memory[1057], memory[1058], memory[1059]};
wire [31:0] memory1060 = {memory[1060], memory[1061], memory[1062], memory[1063]};
wire [31:0] memory1064 = {memory[1064], memory[1065], memory[1066], memory[1067]};
wire [31:0] memory1068 = {memory[1068], memory[1069], memory[1070], memory[1071]};
wire [31:0] memory1072 = {memory[1072], memory[1073], memory[1074], memory[1075]};
wire [31:0] memory1076 = {memory[1076], memory[1077], memory[1078], memory[1079]};
wire [31:0] memory1080 = {memory[1080], memory[1081], memory[1082], memory[1083]};
wire [31:0] memory1084 = {memory[1084], memory[1085], memory[1086], memory[1087]};
wire [31:0] memory1088 = {memory[1088], memory[1089], memory[1090], memory[1091]};
wire [31:0] memory1092 = {memory[1092], memory[1093], memory[1094], memory[1095]};
wire [31:0] memory1096 = {memory[1096], memory[1097], memory[1098], memory[1099]};
wire [31:0] memory1100 = {memory[1100], memory[1101], memory[1102], memory[1103]};
wire [31:0] memory1104 = {memory[1104], memory[1105], memory[1106], memory[1107]};
wire [31:0] memory1108 = {memory[1108], memory[1109], memory[1110], memory[1111]};
wire [31:0] memory1112 = {memory[1112], memory[1113], memory[1114], memory[1115]};
wire [31:0] memory1116 = {memory[1116], memory[1117], memory[1118], memory[1119]};
wire [31:0] memory1120 = {memory[1120], memory[1121], memory[1122], memory[1123]};
wire [31:0] memory1124 = {memory[1124], memory[1125], memory[1126], memory[1127]};
wire [31:0] memory1128 = {memory[1128], memory[1129], memory[1130], memory[1131]};
wire [31:0] memory1132 = {memory[1132], memory[1133], memory[1134], memory[1135]};
wire [31:0] memory1136 = {memory[1136], memory[1137], memory[1138], memory[1139]};
wire [31:0] memory1140 = {memory[1140], memory[1141], memory[1142], memory[1143]};
wire [31:0] memory1144 = {memory[1144], memory[1145], memory[1146], memory[1147]};
wire [31:0] memory1148 = {memory[1148], memory[1149], memory[1150], memory[1151]};
wire [31:0] memory1152 = {memory[1152], memory[1153], memory[1154], memory[1155]};
wire [31:0] memory1156 = {memory[1156], memory[1157], memory[1158], memory[1159]};
wire [31:0] memory1160 = {memory[1160], memory[1161], memory[1162], memory[1163]};
wire [31:0] memory1164 = {memory[1164], memory[1165], memory[1166], memory[1167]};
wire [31:0] memory1168 = {memory[1168], memory[1169], memory[1170], memory[1171]};
wire [31:0] memory1172 = {memory[1172], memory[1173], memory[1174], memory[1175]};
wire [31:0] memory1176 = {memory[1176], memory[1177], memory[1178], memory[1179]};
wire [31:0] memory1180 = {memory[1180], memory[1181], memory[1182], memory[1183]};
wire [31:0] memory1184 = {memory[1184], memory[1185], memory[1186], memory[1187]};
wire [31:0] memory1188 = {memory[1188], memory[1189], memory[1190], memory[1191]};
wire [31:0] memory1192 = {memory[1192], memory[1193], memory[1194], memory[1195]};
wire [31:0] memory1196 = {memory[1196], memory[1197], memory[1198], memory[1199]};
wire [31:0] memory1200 = {memory[1200], memory[1201], memory[1202], memory[1203]};
wire [31:0] memory1204 = {memory[1204], memory[1205], memory[1206], memory[1207]};
wire [31:0] memory1208 = {memory[1208], memory[1209], memory[1210], memory[1211]};
wire [31:0] memory1212 = {memory[1212], memory[1213], memory[1214], memory[1215]};
wire [31:0] memory1216 = {memory[1216], memory[1217], memory[1218], memory[1219]};
wire [31:0] memory1220 = {memory[1220], memory[1221], memory[1222], memory[1223]};
wire [31:0] memory1224 = {memory[1224], memory[1225], memory[1226], memory[1227]};
wire [31:0] memory1228 = {memory[1228], memory[1229], memory[1230], memory[1231]};
wire [31:0] memory1232 = {memory[1232], memory[1233], memory[1234], memory[1235]};
wire [31:0] memory1236 = {memory[1236], memory[1237], memory[1238], memory[1239]};
wire [31:0] memory1240 = {memory[1240], memory[1241], memory[1242], memory[1243]};
wire [31:0] memory1244 = {memory[1244], memory[1245], memory[1246], memory[1247]};
wire [31:0] memory1248 = {memory[1248], memory[1249], memory[1250], memory[1251]};
wire [31:0] memory1252 = {memory[1252], memory[1253], memory[1254], memory[1255]};
wire [31:0] memory1256 = {memory[1256], memory[1257], memory[1258], memory[1259]};
wire [31:0] memory1260 = {memory[1260], memory[1261], memory[1262], memory[1263]};
wire [31:0] memory1264 = {memory[1264], memory[1265], memory[1266], memory[1267]};
wire [31:0] memory1268 = {memory[1268], memory[1269], memory[1270], memory[1271]};
wire [31:0] memory1272 = {memory[1272], memory[1273], memory[1274], memory[1275]};
wire [31:0] memory1276 = {memory[1276], memory[1277], memory[1278], memory[1279]};
wire [31:0] memory1280 = {memory[1280], memory[1281], memory[1282], memory[1283]};
wire [31:0] memory1284 = {memory[1284], memory[1285], memory[1286], memory[1287]};
wire [31:0] memory1288 = {memory[1288], memory[1289], memory[1290], memory[1291]};
wire [31:0] memory1292 = {memory[1292], memory[1293], memory[1294], memory[1295]};
wire [31:0] memory1296 = {memory[1296], memory[1297], memory[1298], memory[1299]};
wire [31:0] memory1300 = {memory[1300], memory[1301], memory[1302], memory[1303]};
wire [31:0] memory1304 = {memory[1304], memory[1305], memory[1306], memory[1307]};
wire [31:0] memory1308 = {memory[1308], memory[1309], memory[1310], memory[1311]};
wire [31:0] memory1312 = {memory[1312], memory[1313], memory[1314], memory[1315]};
wire [31:0] memory1316 = {memory[1316], memory[1317], memory[1318], memory[1319]};
wire [31:0] memory1320 = {memory[1320], memory[1321], memory[1322], memory[1323]};
wire [31:0] memory1324 = {memory[1324], memory[1325], memory[1326], memory[1327]};
wire [31:0] memory1328 = {memory[1328], memory[1329], memory[1330], memory[1331]};
wire [31:0] memory1332 = {memory[1332], memory[1333], memory[1334], memory[1335]};
wire [31:0] memory1336 = {memory[1336], memory[1337], memory[1338], memory[1339]};
wire [31:0] memory1340 = {memory[1340], memory[1341], memory[1342], memory[1343]};
wire [31:0] memory1344 = {memory[1344], memory[1345], memory[1346], memory[1347]};
wire [31:0] memory1348 = {memory[1348], memory[1349], memory[1350], memory[1351]};
wire [31:0] memory1352 = {memory[1352], memory[1353], memory[1354], memory[1355]};
wire [31:0] memory1356 = {memory[1356], memory[1357], memory[1358], memory[1359]};
wire [31:0] memory1360 = {memory[1360], memory[1361], memory[1362], memory[1363]};
wire [31:0] memory1364 = {memory[1364], memory[1365], memory[1366], memory[1367]};
wire [31:0] memory1368 = {memory[1368], memory[1369], memory[1370], memory[1371]};
wire [31:0] memory1372 = {memory[1372], memory[1373], memory[1374], memory[1375]};
wire [31:0] memory1376 = {memory[1376], memory[1377], memory[1378], memory[1379]};
wire [31:0] memory1380 = {memory[1380], memory[1381], memory[1382], memory[1383]};
wire [31:0] memory1384 = {memory[1384], memory[1385], memory[1386], memory[1387]};
wire [31:0] memory1388 = {memory[1388], memory[1389], memory[1390], memory[1391]};
wire [31:0] memory1392 = {memory[1392], memory[1393], memory[1394], memory[1395]};
wire [31:0] memory1396 = {memory[1396], memory[1397], memory[1398], memory[1399]};
wire [31:0] memory1400 = {memory[1400], memory[1401], memory[1402], memory[1403]};
wire [31:0] memory1404 = {memory[1404], memory[1405], memory[1406], memory[1407]};
wire [31:0] memory1408 = {memory[1408], memory[1409], memory[1410], memory[1411]};
wire [31:0] memory1412 = {memory[1412], memory[1413], memory[1414], memory[1415]};
wire [31:0] memory1416 = {memory[1416], memory[1417], memory[1418], memory[1419]};
wire [31:0] memory1420 = {memory[1420], memory[1421], memory[1422], memory[1423]};
wire [31:0] memory1424 = {memory[1424], memory[1425], memory[1426], memory[1427]};
wire [31:0] memory1428 = {memory[1428], memory[1429], memory[1430], memory[1431]};
wire [31:0] memory1432 = {memory[1432], memory[1433], memory[1434], memory[1435]};
wire [31:0] memory1436 = {memory[1436], memory[1437], memory[1438], memory[1439]};
wire [31:0] memory1440 = {memory[1440], memory[1441], memory[1442], memory[1443]};
wire [31:0] memory1444 = {memory[1444], memory[1445], memory[1446], memory[1447]};
wire [31:0] memory1448 = {memory[1448], memory[1449], memory[1450], memory[1451]};
wire [31:0] memory1452 = {memory[1452], memory[1453], memory[1454], memory[1455]};
wire [31:0] memory1456 = {memory[1456], memory[1457], memory[1458], memory[1459]};
wire [31:0] memory1460 = {memory[1460], memory[1461], memory[1462], memory[1463]};
wire [31:0] memory1464 = {memory[1464], memory[1465], memory[1466], memory[1467]};
wire [31:0] memory1468 = {memory[1468], memory[1469], memory[1470], memory[1471]};
wire [31:0] memory1472 = {memory[1472], memory[1473], memory[1474], memory[1475]};
wire [31:0] memory1476 = {memory[1476], memory[1477], memory[1478], memory[1479]};
wire [31:0] memory1480 = {memory[1480], memory[1481], memory[1482], memory[1483]};
wire [31:0] memory1484 = {memory[1484], memory[1485], memory[1486], memory[1487]};
wire [31:0] memory1488 = {memory[1488], memory[1489], memory[1490], memory[1491]};
wire [31:0] memory1492 = {memory[1492], memory[1493], memory[1494], memory[1495]};
wire [31:0] memory1496 = {memory[1496], memory[1497], memory[1498], memory[1499]};
wire [31:0] memory1500 = {memory[1500], memory[1501], memory[1502], memory[1503]};
wire [31:0] memory1504 = {memory[1504], memory[1505], memory[1506], memory[1507]};
wire [31:0] memory1508 = {memory[1508], memory[1509], memory[1510], memory[1511]};
wire [31:0] memory1512 = {memory[1512], memory[1513], memory[1514], memory[1515]};
wire [31:0] memory1516 = {memory[1516], memory[1517], memory[1518], memory[1519]};
wire [31:0] memory1520 = {memory[1520], memory[1521], memory[1522], memory[1523]};
wire [31:0] memory1524 = {memory[1524], memory[1525], memory[1526], memory[1527]};
wire [31:0] memory1528 = {memory[1528], memory[1529], memory[1530], memory[1531]};
wire [31:0] memory1532 = {memory[1532], memory[1533], memory[1534], memory[1535]};
wire [31:0] memory1536 = {memory[1536], memory[1537], memory[1538], memory[1539]};
wire [31:0] memory1540 = {memory[1540], memory[1541], memory[1542], memory[1543]};
wire [31:0] memory1544 = {memory[1544], memory[1545], memory[1546], memory[1547]};
wire [31:0] memory1548 = {memory[1548], memory[1549], memory[1550], memory[1551]};
wire [31:0] memory1552 = {memory[1552], memory[1553], memory[1554], memory[1555]};
wire [31:0] memory1556 = {memory[1556], memory[1557], memory[1558], memory[1559]};
wire [31:0] memory1560 = {memory[1560], memory[1561], memory[1562], memory[1563]};
wire [31:0] memory1564 = {memory[1564], memory[1565], memory[1566], memory[1567]};
wire [31:0] memory1568 = {memory[1568], memory[1569], memory[1570], memory[1571]};
wire [31:0] memory1572 = {memory[1572], memory[1573], memory[1574], memory[1575]};
wire [31:0] memory1576 = {memory[1576], memory[1577], memory[1578], memory[1579]};
wire [31:0] memory1580 = {memory[1580], memory[1581], memory[1582], memory[1583]};
wire [31:0] memory1584 = {memory[1584], memory[1585], memory[1586], memory[1587]};
wire [31:0] memory1588 = {memory[1588], memory[1589], memory[1590], memory[1591]};
wire [31:0] memory1592 = {memory[1592], memory[1593], memory[1594], memory[1595]};
wire [31:0] memory1596 = {memory[1596], memory[1597], memory[1598], memory[1599]};
wire [31:0] memory1600 = {memory[1600], memory[1601], memory[1602], memory[1603]};
wire [31:0] memory1604 = {memory[1604], memory[1605], memory[1606], memory[1607]};
wire [31:0] memory1608 = {memory[1608], memory[1609], memory[1610], memory[1611]};
wire [31:0] memory1612 = {memory[1612], memory[1613], memory[1614], memory[1615]};
wire [31:0] memory1616 = {memory[1616], memory[1617], memory[1618], memory[1619]};
wire [31:0] memory1620 = {memory[1620], memory[1621], memory[1622], memory[1623]};
wire [31:0] memory1624 = {memory[1624], memory[1625], memory[1626], memory[1627]};
wire [31:0] memory1628 = {memory[1628], memory[1629], memory[1630], memory[1631]};
wire [31:0] memory1632 = {memory[1632], memory[1633], memory[1634], memory[1635]};
wire [31:0] memory1636 = {memory[1636], memory[1637], memory[1638], memory[1639]};
wire [31:0] memory1640 = {memory[1640], memory[1641], memory[1642], memory[1643]};
wire [31:0] memory1644 = {memory[1644], memory[1645], memory[1646], memory[1647]};
wire [31:0] memory1648 = {memory[1648], memory[1649], memory[1650], memory[1651]};
wire [31:0] memory1652 = {memory[1652], memory[1653], memory[1654], memory[1655]};
wire [31:0] memory1656 = {memory[1656], memory[1657], memory[1658], memory[1659]};
wire [31:0] memory1660 = {memory[1660], memory[1661], memory[1662], memory[1663]};
wire [31:0] memory1664 = {memory[1664], memory[1665], memory[1666], memory[1667]};
wire [31:0] memory1668 = {memory[1668], memory[1669], memory[1670], memory[1671]};
wire [31:0] memory1672 = {memory[1672], memory[1673], memory[1674], memory[1675]};
wire [31:0] memory1676 = {memory[1676], memory[1677], memory[1678], memory[1679]};
wire [31:0] memory1680 = {memory[1680], memory[1681], memory[1682], memory[1683]};
wire [31:0] memory1684 = {memory[1684], memory[1685], memory[1686], memory[1687]};
wire [31:0] memory1688 = {memory[1688], memory[1689], memory[1690], memory[1691]};
wire [31:0] memory1692 = {memory[1692], memory[1693], memory[1694], memory[1695]};
wire [31:0] memory1696 = {memory[1696], memory[1697], memory[1698], memory[1699]};
wire [31:0] memory1700 = {memory[1700], memory[1701], memory[1702], memory[1703]};
wire [31:0] memory1704 = {memory[1704], memory[1705], memory[1706], memory[1707]};
wire [31:0] memory1708 = {memory[1708], memory[1709], memory[1710], memory[1711]};
wire [31:0] memory1712 = {memory[1712], memory[1713], memory[1714], memory[1715]};
wire [31:0] memory1716 = {memory[1716], memory[1717], memory[1718], memory[1719]};
wire [31:0] memory1720 = {memory[1720], memory[1721], memory[1722], memory[1723]};
wire [31:0] memory1724 = {memory[1724], memory[1725], memory[1726], memory[1727]};
wire [31:0] memory1728 = {memory[1728], memory[1729], memory[1730], memory[1731]};
wire [31:0] memory1732 = {memory[1732], memory[1733], memory[1734], memory[1735]};
wire [31:0] memory1736 = {memory[1736], memory[1737], memory[1738], memory[1739]};
wire [31:0] memory1740 = {memory[1740], memory[1741], memory[1742], memory[1743]};
wire [31:0] memory1744 = {memory[1744], memory[1745], memory[1746], memory[1747]};
wire [31:0] memory1748 = {memory[1748], memory[1749], memory[1750], memory[1751]};
wire [31:0] memory1752 = {memory[1752], memory[1753], memory[1754], memory[1755]};
wire [31:0] memory1756 = {memory[1756], memory[1757], memory[1758], memory[1759]};
wire [31:0] memory1760 = {memory[1760], memory[1761], memory[1762], memory[1763]};
wire [31:0] memory1764 = {memory[1764], memory[1765], memory[1766], memory[1767]};
wire [31:0] memory1768 = {memory[1768], memory[1769], memory[1770], memory[1771]};
wire [31:0] memory1772 = {memory[1772], memory[1773], memory[1774], memory[1775]};
wire [31:0] memory1776 = {memory[1776], memory[1777], memory[1778], memory[1779]};
wire [31:0] memory1780 = {memory[1780], memory[1781], memory[1782], memory[1783]};
wire [31:0] memory1784 = {memory[1784], memory[1785], memory[1786], memory[1787]};
wire [31:0] memory1788 = {memory[1788], memory[1789], memory[1790], memory[1791]};
wire [31:0] memory1792 = {memory[1792], memory[1793], memory[1794], memory[1795]};
wire [31:0] memory1796 = {memory[1796], memory[1797], memory[1798], memory[1799]};
wire [31:0] memory1800 = {memory[1800], memory[1801], memory[1802], memory[1803]};
wire [31:0] memory1804 = {memory[1804], memory[1805], memory[1806], memory[1807]};
wire [31:0] memory1808 = {memory[1808], memory[1809], memory[1810], memory[1811]};
wire [31:0] memory1812 = {memory[1812], memory[1813], memory[1814], memory[1815]};
wire [31:0] memory1816 = {memory[1816], memory[1817], memory[1818], memory[1819]};
wire [31:0] memory1820 = {memory[1820], memory[1821], memory[1822], memory[1823]};
wire [31:0] memory1824 = {memory[1824], memory[1825], memory[1826], memory[1827]};
wire [31:0] memory1828 = {memory[1828], memory[1829], memory[1830], memory[1831]};
wire [31:0] memory1832 = {memory[1832], memory[1833], memory[1834], memory[1835]};
wire [31:0] memory1836 = {memory[1836], memory[1837], memory[1838], memory[1839]};
wire [31:0] memory1840 = {memory[1840], memory[1841], memory[1842], memory[1843]};
wire [31:0] memory1844 = {memory[1844], memory[1845], memory[1846], memory[1847]};
wire [31:0] memory1848 = {memory[1848], memory[1849], memory[1850], memory[1851]};
wire [31:0] memory1852 = {memory[1852], memory[1853], memory[1854], memory[1855]};
wire [31:0] memory1856 = {memory[1856], memory[1857], memory[1858], memory[1859]};
wire [31:0] memory1860 = {memory[1860], memory[1861], memory[1862], memory[1863]};
wire [31:0] memory1864 = {memory[1864], memory[1865], memory[1866], memory[1867]};
wire [31:0] memory1868 = {memory[1868], memory[1869], memory[1870], memory[1871]};
wire [31:0] memory1872 = {memory[1872], memory[1873], memory[1874], memory[1875]};
wire [31:0] memory1876 = {memory[1876], memory[1877], memory[1878], memory[1879]};
wire [31:0] memory1880 = {memory[1880], memory[1881], memory[1882], memory[1883]};
wire [31:0] memory1884 = {memory[1884], memory[1885], memory[1886], memory[1887]};
wire [31:0] memory1888 = {memory[1888], memory[1889], memory[1890], memory[1891]};
wire [31:0] memory1892 = {memory[1892], memory[1893], memory[1894], memory[1895]};
wire [31:0] memory1896 = {memory[1896], memory[1897], memory[1898], memory[1899]};
wire [31:0] memory1900 = {memory[1900], memory[1901], memory[1902], memory[1903]};
wire [31:0] memory1904 = {memory[1904], memory[1905], memory[1906], memory[1907]};
wire [31:0] memory1908 = {memory[1908], memory[1909], memory[1910], memory[1911]};
wire [31:0] memory1912 = {memory[1912], memory[1913], memory[1914], memory[1915]};
wire [31:0] memory1916 = {memory[1916], memory[1917], memory[1918], memory[1919]};
wire [31:0] memory1920 = {memory[1920], memory[1921], memory[1922], memory[1923]};
wire [31:0] memory1924 = {memory[1924], memory[1925], memory[1926], memory[1927]};
wire [31:0] memory1928 = {memory[1928], memory[1929], memory[1930], memory[1931]};
wire [31:0] memory1932 = {memory[1932], memory[1933], memory[1934], memory[1935]};
wire [31:0] memory1936 = {memory[1936], memory[1937], memory[1938], memory[1939]};
wire [31:0] memory1940 = {memory[1940], memory[1941], memory[1942], memory[1943]};
wire [31:0] memory1944 = {memory[1944], memory[1945], memory[1946], memory[1947]};
wire [31:0] memory1948 = {memory[1948], memory[1949], memory[1950], memory[1951]};
wire [31:0] memory1952 = {memory[1952], memory[1953], memory[1954], memory[1955]};
wire [31:0] memory1956 = {memory[1956], memory[1957], memory[1958], memory[1959]};
wire [31:0] memory1960 = {memory[1960], memory[1961], memory[1962], memory[1963]};
wire [31:0] memory1964 = {memory[1964], memory[1965], memory[1966], memory[1967]};
wire [31:0] memory1968 = {memory[1968], memory[1969], memory[1970], memory[1971]};
wire [31:0] memory1972 = {memory[1972], memory[1973], memory[1974], memory[1975]};
wire [31:0] memory1976 = {memory[1976], memory[1977], memory[1978], memory[1979]};
wire [31:0] memory1980 = {memory[1980], memory[1981], memory[1982], memory[1983]};
wire [31:0] memory1984 = {memory[1984], memory[1985], memory[1986], memory[1987]};
wire [31:0] memory1988 = {memory[1988], memory[1989], memory[1990], memory[1991]};
wire [31:0] memory1992 = {memory[1992], memory[1993], memory[1994], memory[1995]};
wire [31:0] memory1996 = {memory[1996], memory[1997], memory[1998], memory[1999]};
wire [31:0] memory2000 = {memory[2000], memory[2001], memory[2002], memory[2003]};
wire [31:0] memory2004 = {memory[2004], memory[2005], memory[2006], memory[2007]};
wire [31:0] memory2008 = {memory[2008], memory[2009], memory[2010], memory[2011]};
wire [31:0] memory2012 = {memory[2012], memory[2013], memory[2014], memory[2015]};
wire [31:0] memory2016 = {memory[2016], memory[2017], memory[2018], memory[2019]};
wire [31:0] memory2020 = {memory[2020], memory[2021], memory[2022], memory[2023]};
wire [31:0] memory2024 = {memory[2024], memory[2025], memory[2026], memory[2027]};
wire [31:0] memory2028 = {memory[2028], memory[2029], memory[2030], memory[2031]};
wire [31:0] memory2032 = {memory[2032], memory[2033], memory[2034], memory[2035]};
wire [31:0] memory2036 = {memory[2036], memory[2037], memory[2038], memory[2039]};
wire [31:0] memory2040 = {memory[2040], memory[2041], memory[2042], memory[2043]};
wire [31:0] memory2044 = {memory[2044], memory[2045], memory[2046], memory[2047]};
wire [31:0] memory2048 = {memory[2048], memory[2049], memory[2050], memory[2051]};
wire [31:0] memory2052 = {memory[2052], memory[2053], memory[2054], memory[2055]};
wire [31:0] memory2056 = {memory[2056], memory[2057], memory[2058], memory[2059]};
wire [31:0] memory2060 = {memory[2060], memory[2061], memory[2062], memory[2063]};
wire [31:0] memory2064 = {memory[2064], memory[2065], memory[2066], memory[2067]};
wire [31:0] memory2068 = {memory[2068], memory[2069], memory[2070], memory[2071]};
wire [31:0] memory2072 = {memory[2072], memory[2073], memory[2074], memory[2075]};
wire [31:0] memory2076 = {memory[2076], memory[2077], memory[2078], memory[2079]};
wire [31:0] memory2080 = {memory[2080], memory[2081], memory[2082], memory[2083]};
wire [31:0] memory2084 = {memory[2084], memory[2085], memory[2086], memory[2087]};
wire [31:0] memory2088 = {memory[2088], memory[2089], memory[2090], memory[2091]};
wire [31:0] memory2092 = {memory[2092], memory[2093], memory[2094], memory[2095]};
wire [31:0] memory2096 = {memory[2096], memory[2097], memory[2098], memory[2099]};
wire [31:0] memory2100 = {memory[2100], memory[2101], memory[2102], memory[2103]};
wire [31:0] memory2104 = {memory[2104], memory[2105], memory[2106], memory[2107]};
wire [31:0] memory2108 = {memory[2108], memory[2109], memory[2110], memory[2111]};
wire [31:0] memory2112 = {memory[2112], memory[2113], memory[2114], memory[2115]};
wire [31:0] memory2116 = {memory[2116], memory[2117], memory[2118], memory[2119]};
wire [31:0] memory2120 = {memory[2120], memory[2121], memory[2122], memory[2123]};
wire [31:0] memory2124 = {memory[2124], memory[2125], memory[2126], memory[2127]};
wire [31:0] memory2128 = {memory[2128], memory[2129], memory[2130], memory[2131]};
wire [31:0] memory2132 = {memory[2132], memory[2133], memory[2134], memory[2135]};
wire [31:0] memory2136 = {memory[2136], memory[2137], memory[2138], memory[2139]};
wire [31:0] memory2140 = {memory[2140], memory[2141], memory[2142], memory[2143]};
wire [31:0] memory2144 = {memory[2144], memory[2145], memory[2146], memory[2147]};
wire [31:0] memory2148 = {memory[2148], memory[2149], memory[2150], memory[2151]};
wire [31:0] memory2152 = {memory[2152], memory[2153], memory[2154], memory[2155]};
wire [31:0] memory2156 = {memory[2156], memory[2157], memory[2158], memory[2159]};
wire [31:0] memory2160 = {memory[2160], memory[2161], memory[2162], memory[2163]};
wire [31:0] memory2164 = {memory[2164], memory[2165], memory[2166], memory[2167]};
wire [31:0] memory2168 = {memory[2168], memory[2169], memory[2170], memory[2171]};
wire [31:0] memory2172 = {memory[2172], memory[2173], memory[2174], memory[2175]};
wire [31:0] memory2176 = {memory[2176], memory[2177], memory[2178], memory[2179]};
wire [31:0] memory2180 = {memory[2180], memory[2181], memory[2182], memory[2183]};
wire [31:0] memory2184 = {memory[2184], memory[2185], memory[2186], memory[2187]};
wire [31:0] memory2188 = {memory[2188], memory[2189], memory[2190], memory[2191]};
wire [31:0] memory2192 = {memory[2192], memory[2193], memory[2194], memory[2195]};
wire [31:0] memory2196 = {memory[2196], memory[2197], memory[2198], memory[2199]};
wire [31:0] memory2200 = {memory[2200], memory[2201], memory[2202], memory[2203]};
wire [31:0] memory2204 = {memory[2204], memory[2205], memory[2206], memory[2207]};
wire [31:0] memory2208 = {memory[2208], memory[2209], memory[2210], memory[2211]};
wire [31:0] memory2212 = {memory[2212], memory[2213], memory[2214], memory[2215]};
wire [31:0] memory2216 = {memory[2216], memory[2217], memory[2218], memory[2219]};
wire [31:0] memory2220 = {memory[2220], memory[2221], memory[2222], memory[2223]};
wire [31:0] memory2224 = {memory[2224], memory[2225], memory[2226], memory[2227]};
wire [31:0] memory2228 = {memory[2228], memory[2229], memory[2230], memory[2231]};
wire [31:0] memory2232 = {memory[2232], memory[2233], memory[2234], memory[2235]};
wire [31:0] memory2236 = {memory[2236], memory[2237], memory[2238], memory[2239]};
wire [31:0] memory2240 = {memory[2240], memory[2241], memory[2242], memory[2243]};
wire [31:0] memory2244 = {memory[2244], memory[2245], memory[2246], memory[2247]};
wire [31:0] memory2248 = {memory[2248], memory[2249], memory[2250], memory[2251]};
wire [31:0] memory2252 = {memory[2252], memory[2253], memory[2254], memory[2255]};
wire [31:0] memory2256 = {memory[2256], memory[2257], memory[2258], memory[2259]};
wire [31:0] memory2260 = {memory[2260], memory[2261], memory[2262], memory[2263]};
wire [31:0] memory2264 = {memory[2264], memory[2265], memory[2266], memory[2267]};
wire [31:0] memory2268 = {memory[2268], memory[2269], memory[2270], memory[2271]};
wire [31:0] memory2272 = {memory[2272], memory[2273], memory[2274], memory[2275]};
wire [31:0] memory2276 = {memory[2276], memory[2277], memory[2278], memory[2279]};
// Ponte para debug da memória dat[0] até dat[1023], agrupando em words de 32 bits
wire [31:0] memory25996 = {memory[25996], memory[25997], memory[25998], memory[25999]};
wire [31:0] memory26000 = {memory[26000], memory[26001], memory[26002], memory[26003]};
wire [31:0] memory26004 = {memory[26004], memory[26005], memory[26006], memory[26007]};
wire [31:0] memory26008 = {memory[26008], memory[26009], memory[26010], memory[26011]};
wire [31:0] memory26012 = {memory[26012], memory[26013], memory[26014], memory[26015]};
wire [31:0] memory26016 = {memory[26016], memory[26017], memory[26018], memory[26019]};
wire [31:0] memory26020 = {memory[26020], memory[26021], memory[26022], memory[26023]};
wire [31:0] memory26024 = {memory[26024], memory[26025], memory[26026], memory[26027]};
wire [31:0] memory26028 = {memory[26028], memory[26029], memory[26030], memory[26031]};
wire [31:0] memory26032 = {memory[26032], memory[26033], memory[26034], memory[26035]};
wire [31:0] memory26036 = {memory[26036], memory[26037], memory[26038], memory[26039]};
wire [31:0] memory26040 = {memory[26040], memory[26041], memory[26042], memory[26043]};
wire [31:0] memory26044 = {memory[26044], memory[26045], memory[26046], memory[26047]};
wire [31:0] memory26048 = {memory[26048], memory[26049], memory[26050], memory[26051]};
wire [31:0] memory26052 = {memory[26052], memory[26053], memory[26054], memory[26055]};
wire [31:0] memory26056 = {memory[26056], memory[26057], memory[26058], memory[26059]};
wire [31:0] memory26060 = {memory[26060], memory[26061], memory[26062], memory[26063]};
wire [31:0] memory26064 = {memory[26064], memory[26065], memory[26066], memory[26067]};
wire [31:0] memory26068 = {memory[26068], memory[26069], memory[26070], memory[26071]};
wire [31:0] memory26072 = {memory[26072], memory[26073], memory[26074], memory[26075]};
wire [31:0] memory26076 = {memory[26076], memory[26077], memory[26078], memory[26079]};
wire [31:0] memory26080 = {memory[26080], memory[26081], memory[26082], memory[26083]};
wire [31:0] memory26084 = {memory[26084], memory[26085], memory[26086], memory[26087]};
wire [31:0] memory26088 = {memory[26088], memory[26089], memory[26090], memory[26091]};
wire [31:0] memory26092 = {memory[26092], memory[26093], memory[26094], memory[26095]};
wire [31:0] memory26096 = {memory[26096], memory[26097], memory[26098], memory[26099]};
wire [31:0] memory26100 = {memory[26100], memory[26101], memory[26102], memory[26103]};
wire [31:0] memory26104 = {memory[26104], memory[26105], memory[26106], memory[26107]};
wire [31:0] memory26108 = {memory[26108], memory[26109], memory[26110], memory[26111]};
wire [31:0] memory26112 = {memory[26112], memory[26113], memory[26114], memory[26115]};
wire [31:0] memory26116 = {memory[26116], memory[26117], memory[26118], memory[26119]};
wire [31:0] memory26120 = {memory[26120], memory[26121], memory[26122], memory[26123]};
wire [31:0] memory26124 = {memory[26124], memory[26125], memory[26126], memory[26127]};
wire [31:0] memory26128 = {memory[26128], memory[26129], memory[26130], memory[26131]};
wire [31:0] memory26132 = {memory[26132], memory[26133], memory[26134], memory[26135]};
wire [31:0] memory26136 = {memory[26136], memory[26137], memory[26138], memory[26139]};
wire [31:0] memory26140 = {memory[26140], memory[26141], memory[26142], memory[26143]};
wire [31:0] memory26144 = {memory[26144], memory[26145], memory[26146], memory[26147]};
wire [31:0] memory26148 = {memory[26148], memory[26149], memory[26150], memory[26151]};
wire [31:0] memory26152 = {memory[26152], memory[26153], memory[26154], memory[26155]};
wire [31:0] memory26156 = {memory[26156], memory[26157], memory[26158], memory[26159]};
wire [31:0] memory26160 = {memory[26160], memory[26161], memory[26162], memory[26163]};
wire [31:0] memory26164 = {memory[26164], memory[26165], memory[26166], memory[26167]};
wire [31:0] memory26168 = {memory[26168], memory[26169], memory[26170], memory[26171]};
wire [31:0] memory26172 = {memory[26172], memory[26173], memory[26174], memory[26175]};
wire [31:0] memory26176 = {memory[26176], memory[26177], memory[26178], memory[26179]};
wire [31:0] memory26180 = {memory[26180], memory[26181], memory[26182], memory[26183]};
wire [31:0] memory26184 = {memory[26184], memory[26185], memory[26186], memory[26187]};
wire [31:0] memory26188 = {memory[26188], memory[26189], memory[26190], memory[26191]};
wire [31:0] memory26192 = {memory[26192], memory[26193], memory[26194], memory[26195]};
wire [31:0] memory26196 = {memory[26196], memory[26197], memory[26198], memory[26199]};
wire [31:0] memory26200 = {memory[26200], memory[26201], memory[26202], memory[26203]};
wire [31:0] memory26204 = {memory[26204], memory[26205], memory[26206], memory[26207]};
wire [31:0] memory26208 = {memory[26208], memory[26209], memory[26210], memory[26211]};
wire [31:0] memory26212 = {memory[26212], memory[26213], memory[26214], memory[26215]};
wire [31:0] memory26216 = {memory[26216], memory[26217], memory[26218], memory[26219]};
wire [31:0] memory26220 = {memory[26220], memory[26221], memory[26222], memory[26223]};
wire [31:0] memory26224 = {memory[26224], memory[26225], memory[26226], memory[26227]};
wire [31:0] memory26228 = {memory[26228], memory[26229], memory[26230], memory[26231]};
wire [31:0] memory26232 = {memory[26232], memory[26233], memory[26234], memory[26235]};
wire [31:0] memory26236 = {memory[26236], memory[26237], memory[26238], memory[26239]};
wire [31:0] memory26240 = {memory[26240], memory[26241], memory[26242], memory[26243]};
wire [31:0] memory26244 = {memory[26244], memory[26245], memory[26246], memory[26247]};
wire [31:0] memory26248 = {memory[26248], memory[26249], memory[26250], memory[26251]};
wire [31:0] memory26252 = {memory[26252], memory[26253], memory[26254], memory[26255]};
wire [31:0] memory26256 = {memory[26256], memory[26257], memory[26258], memory[26259]};
wire [31:0] memory26260 = {memory[26260], memory[26261], memory[26262], memory[26263]};
wire [31:0] memory26264 = {memory[26264], memory[26265], memory[26266], memory[26267]};
wire [31:0] memory26268 = {memory[26268], memory[26269], memory[26270], memory[26271]};
wire [31:0] memory26272 = {memory[26272], memory[26273], memory[26274], memory[26275]};
wire [31:0] memory26276 = {memory[26276], memory[26277], memory[26278], memory[26279]};
wire [31:0] memory26280 = {memory[26280], memory[26281], memory[26282], memory[26283]};
wire [31:0] memory26284 = {memory[26284], memory[26285], memory[26286], memory[26287]};
wire [31:0] memory26288 = {memory[26288], memory[26289], memory[26290], memory[26291]};
wire [31:0] memory26292 = {memory[26292], memory[26293], memory[26294], memory[26295]};
wire [31:0] memory26296 = {memory[26296], memory[26297], memory[26298], memory[26299]};
wire [31:0] memory26300 = {memory[26300], memory[26301], memory[26302], memory[26303]};
wire [31:0] memory26304 = {memory[26304], memory[26305], memory[26306], memory[26307]};
wire [31:0] memory26308 = {memory[26308], memory[26309], memory[26310], memory[26311]};
wire [31:0] memory26312 = {memory[26312], memory[26313], memory[26314], memory[26315]};
wire [31:0] memory26316 = {memory[26316], memory[26317], memory[26318], memory[26319]};
wire [31:0] memory26320 = {memory[26320], memory[26321], memory[26322], memory[26323]};
wire [31:0] memory26324 = {memory[26324], memory[26325], memory[26326], memory[26327]};
wire [31:0] memory26328 = {memory[26328], memory[26329], memory[26330], memory[26331]};
wire [31:0] memory26332 = {memory[26332], memory[26333], memory[26334], memory[26335]};
wire [31:0] memory26336 = {memory[26336], memory[26337], memory[26338], memory[26339]};
wire [31:0] memory26340 = {memory[26340], memory[26341], memory[26342], memory[26343]};
wire [31:0] memory26344 = {memory[26344], memory[26345], memory[26346], memory[26347]};
wire [31:0] memory26348 = {memory[26348], memory[26349], memory[26350], memory[26351]};
wire [31:0] memory26352 = {memory[26352], memory[26353], memory[26354], memory[26355]};
wire [31:0] memory26356 = {memory[26356], memory[26357], memory[26358], memory[26359]};
wire [31:0] memory26360 = {memory[26360], memory[26361], memory[26362], memory[26363]};
wire [31:0] memory26364 = {memory[26364], memory[26365], memory[26366], memory[26367]};
wire [31:0] memory26368 = {memory[26368], memory[26369], memory[26370], memory[26371]};
wire [31:0] memory26372 = {memory[26372], memory[26373], memory[26374], memory[26375]};
wire [31:0] memory26376 = {memory[26376], memory[26377], memory[26378], memory[26379]};
wire [31:0] memory26380 = {memory[26380], memory[26381], memory[26382], memory[26383]};
wire [31:0] memory26384 = {memory[26384], memory[26385], memory[26386], memory[26387]};
wire [31:0] memory26388 = {memory[26388], memory[26389], memory[26390], memory[26391]};
wire [31:0] memory26392 = {memory[26392], memory[26393], memory[26394], memory[26395]};
wire [31:0] memory26396 = {memory[26396], memory[26397], memory[26398], memory[26399]};
wire [31:0] memory26400 = {memory[26400], memory[26401], memory[26402], memory[26403]};
wire [31:0] memory26404 = {memory[26404], memory[26405], memory[26406], memory[26407]};
wire [31:0] memory26408 = {memory[26408], memory[26409], memory[26410], memory[26411]};
wire [31:0] memory26412 = {memory[26412], memory[26413], memory[26414], memory[26415]};
wire [31:0] memory26416 = {memory[26416], memory[26417], memory[26418], memory[26419]};
wire [31:0] memory26420 = {memory[26420], memory[26421], memory[26422], memory[26423]};
wire [31:0] memory26424 = {memory[26424], memory[26425], memory[26426], memory[26427]};
wire [31:0] memory26428 = {memory[26428], memory[26429], memory[26430], memory[26431]};
wire [31:0] memory26432 = {memory[26432], memory[26433], memory[26434], memory[26435]};
wire [31:0] memory26436 = {memory[26436], memory[26437], memory[26438], memory[26439]};
wire [31:0] memory26440 = {memory[26440], memory[26441], memory[26442], memory[26443]};
wire [31:0] memory26444 = {memory[26444], memory[26445], memory[26446], memory[26447]};
wire [31:0] memory26448 = {memory[26448], memory[26449], memory[26450], memory[26451]};
wire [31:0] memory26452 = {memory[26452], memory[26453], memory[26454], memory[26455]};
wire [31:0] memory26456 = {memory[26456], memory[26457], memory[26458], memory[26459]};
wire [31:0] memory26460 = {memory[26460], memory[26461], memory[26462], memory[26463]};
wire [31:0] memory26464 = {memory[26464], memory[26465], memory[26466], memory[26467]};
wire [31:0] memory26468 = {memory[26468], memory[26469], memory[26470], memory[26471]};
wire [31:0] memory26472 = {memory[26472], memory[26473], memory[26474], memory[26475]};
wire [31:0] memory26476 = {memory[26476], memory[26477], memory[26478], memory[26479]};
wire [31:0] memory26480 = {memory[26480], memory[26481], memory[26482], memory[26483]};
wire [31:0] memory26484 = {memory[26484], memory[26485], memory[26486], memory[26487]};
wire [31:0] memory26488 = {memory[26488], memory[26489], memory[26490], memory[26491]};
wire [31:0] memory26492 = {memory[26492], memory[26493], memory[26494], memory[26495]};
wire [31:0] memory26496 = {memory[26496], memory[26497], memory[26498], memory[26499]};
wire [31:0] memory26500 = {memory[26500], memory[26501], memory[26502], memory[26503]};
wire [31:0] memory26504 = {memory[26504], memory[26505], memory[26506], memory[26507]};
wire [31:0] memory26508 = {memory[26508], memory[26509], memory[26510], memory[26511]};
wire [31:0] memory26512 = {memory[26512], memory[26513], memory[26514], memory[26515]};
wire [31:0] memory26516 = {memory[26516], memory[26517], memory[26518], memory[26519]};
wire [31:0] memory26520 = {memory[26520], memory[26521], memory[26522], memory[26523]};
wire [31:0] memory26524 = {memory[26524], memory[26525], memory[26526], memory[26527]};
wire [31:0] memory26528 = {memory[26528], memory[26529], memory[26530], memory[26531]};
wire [31:0] memory26532 = {memory[26532], memory[26533], memory[26534], memory[26535]};
wire [31:0] memory26536 = {memory[26536], memory[26537], memory[26538], memory[26539]};
wire [31:0] memory26540 = {memory[26540], memory[26541], memory[26542], memory[26543]};
wire [31:0] memory26544 = {memory[26544], memory[26545], memory[26546], memory[26547]};
wire [31:0] memory26548 = {memory[26548], memory[26549], memory[26550], memory[26551]};
wire [31:0] memory26552 = {memory[26552], memory[26553], memory[26554], memory[26555]};
wire [31:0] memory26556 = {memory[26556], memory[26557], memory[26558], memory[26559]};
wire [31:0] memory26560 = {memory[26560], memory[26561], memory[26562], memory[26563]};
wire [31:0] memory26564 = {memory[26564], memory[26565], memory[26566], memory[26567]};
wire [31:0] memory26568 = {memory[26568], memory[26569], memory[26570], memory[26571]};
wire [31:0] memory26572 = {memory[26572], memory[26573], memory[26574], memory[26575]};
wire [31:0] memory26576 = {memory[26576], memory[26577], memory[26578], memory[26579]};
wire [31:0] memory26580 = {memory[26580], memory[26581], memory[26582], memory[26583]};
wire [31:0] memory26584 = {memory[26584], memory[26585], memory[26586], memory[26587]};
wire [31:0] memory26588 = {memory[26588], memory[26589], memory[26590], memory[26591]};
wire [31:0] memory26592 = {memory[26592], memory[26593], memory[26594], memory[26595]};
wire [31:0] memory26596 = {memory[26596], memory[26597], memory[26598], memory[26599]};
wire [31:0] memory26600 = {memory[26600], memory[26601], memory[26602], memory[26603]};
wire [31:0] memory26604 = {memory[26604], memory[26605], memory[26606], memory[26607]};
wire [31:0] memory26608 = {memory[26608], memory[26609], memory[26610], memory[26611]};
wire [31:0] memory26612 = {memory[26612], memory[26613], memory[26614], memory[26615]};
wire [31:0] memory26616 = {memory[26616], memory[26617], memory[26618], memory[26619]};
wire [31:0] memory26620 = {memory[26620], memory[26621], memory[26622], memory[26623]};
wire [31:0] memory26624 = {memory[26624], memory[26625], memory[26626], memory[26627]};
wire [31:0] memory26628 = {memory[26628], memory[26629], memory[26630], memory[26631]};
wire [31:0] memory26632 = {memory[26632], memory[26633], memory[26634], memory[26635]};
wire [31:0] memory26636 = {memory[26636], memory[26637], memory[26638], memory[26639]};
wire [31:0] memory26640 = {memory[26640], memory[26641], memory[26642], memory[26643]};
wire [31:0] memory26644 = {memory[26644], memory[26645], memory[26646], memory[26647]};
wire [31:0] memory26648 = {memory[26648], memory[26649], memory[26650], memory[26651]};
wire [31:0] memory26652 = {memory[26652], memory[26653], memory[26654], memory[26655]};
wire [31:0] memory26656 = {memory[26656], memory[26657], memory[26658], memory[26659]};
wire [31:0] memory26660 = {memory[26660], memory[26661], memory[26662], memory[26663]};
wire [31:0] memory26664 = {memory[26664], memory[26665], memory[26666], memory[26667]};
wire [31:0] memory26668 = {memory[26668], memory[26669], memory[26670], memory[26671]};
wire [31:0] memory26672 = {memory[26672], memory[26673], memory[26674], memory[26675]};
wire [31:0] memory26676 = {memory[26676], memory[26677], memory[26678], memory[26679]};
wire [31:0] memory26680 = {memory[26680], memory[26681], memory[26682], memory[26683]};
wire [31:0] memory26684 = {memory[26684], memory[26685], memory[26686], memory[26687]};
wire [31:0] memory26688 = {memory[26688], memory[26689], memory[26690], memory[26691]};
wire [31:0] memory26692 = {memory[26692], memory[26693], memory[26694], memory[26695]};
wire [31:0] memory26696 = {memory[26696], memory[26697], memory[26698], memory[26699]};
wire [31:0] memory26700 = {memory[26700], memory[26701], memory[26702], memory[26703]};
wire [31:0] memory26704 = {memory[26704], memory[26705], memory[26706], memory[26707]};
wire [31:0] memory26708 = {memory[26708], memory[26709], memory[26710], memory[26711]};
wire [31:0] memory26712 = {memory[26712], memory[26713], memory[26714], memory[26715]};
wire [31:0] memory26716 = {memory[26716], memory[26717], memory[26718], memory[26719]};
wire [31:0] memory26720 = {memory[26720], memory[26721], memory[26722], memory[26723]};
wire [31:0] memory26724 = {memory[26724], memory[26725], memory[26726], memory[26727]};
wire [31:0] memory26728 = {memory[26728], memory[26729], memory[26730], memory[26731]};
wire [31:0] memory26732 = {memory[26732], memory[26733], memory[26734], memory[26735]};
wire [31:0] memory26736 = {memory[26736], memory[26737], memory[26738], memory[26739]};
wire [31:0] memory26740 = {memory[26740], memory[26741], memory[26742], memory[26743]};
wire [31:0] memory26744 = {memory[26744], memory[26745], memory[26746], memory[26747]};
wire [31:0] memory26748 = {memory[26748], memory[26749], memory[26750], memory[26751]};
wire [31:0] memory26752 = {memory[26752], memory[26753], memory[26754], memory[26755]};
wire [31:0] memory26756 = {memory[26756], memory[26757], memory[26758], memory[26759]};
wire [31:0] memory26760 = {memory[26760], memory[26761], memory[26762], memory[26763]};
wire [31:0] memory26764 = {memory[26764], memory[26765], memory[26766], memory[26767]};
wire [31:0] memory26768 = {memory[26768], memory[26769], memory[26770], memory[26771]};
wire [31:0] memory26772 = {memory[26772], memory[26773], memory[26774], memory[26775]};
wire [31:0] memory26776 = {memory[26776], memory[26777], memory[26778], memory[26779]};
wire [31:0] memory26780 = {memory[26780], memory[26781], memory[26782], memory[26783]};
wire [31:0] memory26784 = {memory[26784], memory[26785], memory[26786], memory[26787]};
wire [31:0] memory26788 = {memory[26788], memory[26789], memory[26790], memory[26791]};
wire [31:0] memory26792 = {memory[26792], memory[26793], memory[26794], memory[26795]};
wire [31:0] memory26796 = {memory[26796], memory[26797], memory[26798], memory[26799]};
wire [31:0] memory26800 = {memory[26800], memory[26801], memory[26802], memory[26803]};
wire [31:0] memory26804 = {memory[26804], memory[26805], memory[26806], memory[26807]};
wire [31:0] memory26808 = {memory[26808], memory[26809], memory[26810], memory[26811]};
wire [31:0] memory26812 = {memory[26812], memory[26813], memory[26814], memory[26815]};
wire [31:0] memory26816 = {memory[26816], memory[26817], memory[26818], memory[26819]};
wire [31:0] memory26820 = {memory[26820], memory[26821], memory[26822], memory[26823]};
wire [31:0] memory26824 = {memory[26824], memory[26825], memory[26826], memory[26827]};
wire [31:0] memory26828 = {memory[26828], memory[26829], memory[26830], memory[26831]};
wire [31:0] memory26832 = {memory[26832], memory[26833], memory[26834], memory[26835]};
wire [31:0] memory26836 = {memory[26836], memory[26837], memory[26838], memory[26839]};
wire [31:0] memory26840 = {memory[26840], memory[26841], memory[26842], memory[26843]};
wire [31:0] memory26844 = {memory[26844], memory[26845], memory[26846], memory[26847]};
wire [31:0] memory26848 = {memory[26848], memory[26849], memory[26850], memory[26851]};
wire [31:0] memory26852 = {memory[26852], memory[26853], memory[26854], memory[26855]};
wire [31:0] memory26856 = {memory[26856], memory[26857], memory[26858], memory[26859]};
wire [31:0] memory26860 = {memory[26860], memory[26861], memory[26862], memory[26863]};
wire [31:0] memory26864 = {memory[26864], memory[26865], memory[26866], memory[26867]};
wire [31:0] memory26868 = {memory[26868], memory[26869], memory[26870], memory[26871]};
wire [31:0] memory26872 = {memory[26872], memory[26873], memory[26874], memory[26875]};
wire [31:0] memory26876 = {memory[26876], memory[26877], memory[26878], memory[26879]};
wire [31:0] memory26880 = {memory[26880], memory[26881], memory[26882], memory[26883]};
wire [31:0] memory26884 = {memory[26884], memory[26885], memory[26886], memory[26887]};
wire [31:0] memory26888 = {memory[26888], memory[26889], memory[26890], memory[26891]};
wire [31:0] memory26892 = {memory[26892], memory[26893], memory[26894], memory[26895]};
wire [31:0] memory26896 = {memory[26896], memory[26897], memory[26898], memory[26899]};
wire [31:0] memory26900 = {memory[26900], memory[26901], memory[26902], memory[26903]};
wire [31:0] memory26904 = {memory[26904], memory[26905], memory[26906], memory[26907]};
wire [31:0] memory26908 = {memory[26908], memory[26909], memory[26910], memory[26911]};
wire [31:0] memory26912 = {memory[26912], memory[26913], memory[26914], memory[26915]};
wire [31:0] memory26916 = {memory[26916], memory[26917], memory[26918], memory[26919]};
wire [31:0] memory26920 = {memory[26920], memory[26921], memory[26922], memory[26923]};
wire [31:0] memory26924 = {memory[26924], memory[26925], memory[26926], memory[26927]};
wire [31:0] memory26928 = {memory[26928], memory[26929], memory[26930], memory[26931]};
wire [31:0] memory26932 = {memory[26932], memory[26933], memory[26934], memory[26935]};
wire [31:0] memory26936 = {memory[26936], memory[26937], memory[26938], memory[26939]};
wire [31:0] memory26940 = {memory[26940], memory[26941], memory[26942], memory[26943]};
wire [31:0] memory26944 = {memory[26944], memory[26945], memory[26946], memory[26947]};
wire [31:0] memory26948 = {memory[26948], memory[26949], memory[26950], memory[26951]};
wire [31:0] memory26952 = {memory[26952], memory[26953], memory[26954], memory[26955]};
wire [31:0] memory26956 = {memory[26956], memory[26957], memory[26958], memory[26959]};
wire [31:0] memory26960 = {memory[26960], memory[26961], memory[26962], memory[26963]};
wire [31:0] memory26964 = {memory[26964], memory[26965], memory[26966], memory[26967]};
wire [31:0] memory26968 = {memory[26968], memory[26969], memory[26970], memory[26971]};
wire [31:0] memory26972 = {memory[26972], memory[26973], memory[26974], memory[26975]};
wire [31:0] memory26976 = {memory[26976], memory[26977], memory[26978], memory[26979]};
wire [31:0] memory26980 = {memory[26980], memory[26981], memory[26982], memory[26983]};
wire [31:0] memory26984 = {memory[26984], memory[26985], memory[26986], memory[26987]};
wire [31:0] memory26988 = {memory[26988], memory[26989], memory[26990], memory[26991]};
wire [31:0] memory26992 = {memory[26992], memory[26993], memory[26994], memory[26995]};
wire [31:0] memory26996 = {memory[26996], memory[26997], memory[26998], memory[26999]};
wire [31:0] memory27000 = {memory[27000], memory[27001], memory[27002], memory[27003]};
wire [31:0] memory27004 = {memory[27004], memory[27005], memory[27006], memory[27007]};
wire [31:0] memory27008 = {memory[27008], memory[27009], memory[27010], memory[27011]};
wire [31:0] memory27012 = {memory[27012], memory[27013], memory[27014], memory[27015]};
wire [31:0] memory27016 = {memory[27016], memory[27017], memory[27018], memory[27019]};
wire [31:0] memory27020 = {memory[27020], memory[27021], memory[27022], memory[27023]};
wire [31:0] memory27024 = {memory[27024], memory[27025], memory[27026], memory[27027]};
wire [31:0] memory27028 = {memory[27028], memory[27029], memory[27030], memory[27031]};
wire [31:0] memory27032 = {memory[27032], memory[27033], memory[27034], memory[27035]};
wire [31:0] memory27036 = {memory[27036], memory[27037], memory[27038], memory[27039]};
wire [31:0] memory27040 = {memory[27040], memory[27041], memory[27042], memory[27043]};
wire [31:0] memory27044 = {memory[27044], memory[27045], memory[27046], memory[27047]};
wire [31:0] memory27048 = {memory[27048], memory[27049], memory[27050], memory[27051]};
wire [31:0] memory27052 = {memory[27052], memory[27053], memory[27054], memory[27055]};
wire [31:0] memory27056 = {memory[27056], memory[27057], memory[27058], memory[27059]};
wire [31:0] memory27060 = {memory[27060], memory[27061], memory[27062], memory[27063]};
wire [31:0] memory27064 = {memory[27064], memory[27065], memory[27066], memory[27067]};
wire [31:0] memory27068 = {memory[27068], memory[27069], memory[27070], memory[27071]};
wire [31:0] memory27072 = {memory[27072], memory[27073], memory[27074], memory[27075]};
wire [31:0] memory27076 = {memory[27076], memory[27077], memory[27078], memory[27079]};
wire [31:0] memory27080 = {memory[27080], memory[27081], memory[27082], memory[27083]};
wire [31:0] memory27084 = {memory[27084], memory[27085], memory[27086], memory[27087]};
wire [31:0] memory27088 = {memory[27088], memory[27089], memory[27090], memory[27091]};
wire [31:0] memory27092 = {memory[27092], memory[27093], memory[27094], memory[27095]};
wire [31:0] memory27096 = {memory[27096], memory[27097], memory[27098], memory[27099]};
wire [31:0] memory27100 = {memory[27100], memory[27101], memory[27102], memory[27103]};
wire [31:0] memory27104 = {memory[27104], memory[27105], memory[27106], memory[27107]};
wire [31:0] memory27108 = {memory[27108], memory[27109], memory[27110], memory[27111]};
wire [31:0] memory27112 = {memory[27112], memory[27113], memory[27114], memory[27115]};
wire [31:0] memory27116 = {memory[27116], memory[27117], memory[27118], memory[27119]};
wire [31:0] memory27120 = {memory[27120], memory[27121], memory[27122], memory[27123]};
wire [31:0] memory27124 = {memory[27124], memory[27125], memory[27126], memory[27127]};
wire [31:0] memory27128 = {memory[27128], memory[27129], memory[27130], memory[27131]};
wire [31:0] memory27132 = {memory[27132], memory[27133], memory[27134], memory[27135]};
wire [31:0] memory27136 = {memory[27136], memory[27137], memory[27138], memory[27139]};
wire [31:0] memory27140 = {memory[27140], memory[27141], memory[27142], memory[27143]};
wire [31:0] memory27144 = {memory[27144], memory[27145], memory[27146], memory[27147]};
wire [31:0] memory27148 = {memory[27148], memory[27149], memory[27150], memory[27151]};
wire [31:0] memory27152 = {memory[27152], memory[27153], memory[27154], memory[27155]};
wire [31:0] memory27156 = {memory[27156], memory[27157], memory[27158], memory[27159]};
wire [31:0] memory27160 = {memory[27160], memory[27161], memory[27162], memory[27163]};
wire [31:0] memory27164 = {memory[27164], memory[27165], memory[27166], memory[27167]};
wire [31:0] memory27168 = {memory[27168], memory[27169], memory[27170], memory[27171]};
wire [31:0] memory27172 = {memory[27172], memory[27173], memory[27174], memory[27175]};
wire [31:0] memory27176 = {memory[27176], memory[27177], memory[27178], memory[27179]};
wire [31:0] memory27180 = {memory[27180], memory[27181], memory[27182], memory[27183]};
wire [31:0] memory27184 = {memory[27184], memory[27185], memory[27186], memory[27187]};
wire [31:0] memory27188 = {memory[27188], memory[27189], memory[27190], memory[27191]};
wire [31:0] memory27192 = {memory[27192], memory[27193], memory[27194], memory[27195]};
wire [31:0] memory27196 = {memory[27196], memory[27197], memory[27198], memory[27199]};
wire [31:0] memory27200 = {memory[27200], memory[27201], memory[27202], memory[27203]};
wire [31:0] memory27204 = {memory[27204], memory[27205], memory[27206], memory[27207]};
wire [31:0] memory27208 = {memory[27208], memory[27209], memory[27210], memory[27211]};
wire [31:0] memory27212 = {memory[27212], memory[27213], memory[27214], memory[27215]};
wire [31:0] memory27216 = {memory[27216], memory[27217], memory[27218], memory[27219]};
wire [31:0] memory27220 = {memory[27220], memory[27221], memory[27222], memory[27223]};
wire [31:0] memory27224 = {memory[27224], memory[27225], memory[27226], memory[27227]};
wire [31:0] memory27228 = {memory[27228], memory[27229], memory[27230], memory[27231]};
wire [31:0] memory27232 = {memory[27232], memory[27233], memory[27234], memory[27235]};
wire [31:0] memory27236 = {memory[27236], memory[27237], memory[27238], memory[27239]};
wire [31:0] memory27240 = {memory[27240], memory[27241], memory[27242], memory[27243]};
wire [31:0] memory27244 = {memory[27244], memory[27245], memory[27246], memory[27247]};
wire [31:0] memory27248 = {memory[27248], memory[27249], memory[27250], memory[27251]};
wire [31:0] memory27252 = {memory[27252], memory[27253], memory[27254], memory[27255]};
wire [31:0] memory27256 = {memory[27256], memory[27257], memory[27258], memory[27259]};
wire [31:0] memory27260 = {memory[27260], memory[27261], memory[27262], memory[27263]};
wire [31:0] memory27264 = {memory[27264], memory[27265], memory[27266], memory[27267]};
wire [31:0] memory27268 = {memory[27268], memory[27269], memory[27270], memory[27271]};
wire [31:0] memory27272 = {memory[27272], memory[27273], memory[27274], memory[27275]};
wire [31:0] memory27276 = {memory[27276], memory[27277], memory[27278], memory[27279]};
wire [31:0] memory27280 = {memory[27280], memory[27281], memory[27282], memory[27283]};
wire [31:0] memory27284 = {memory[27284], memory[27285], memory[27286], memory[27287]};
wire [31:0] memory27288 = {memory[27288], memory[27289], memory[27290], memory[27291]};
wire [31:0] memory27292 = {memory[27292], memory[27293], memory[27294], memory[27295]};
wire [31:0] memory27296 = {memory[27296], memory[27297], memory[27298], memory[27299]};
wire [31:0] memory27300 = {memory[27300], memory[27301], memory[27302], memory[27303]};
wire [31:0] memory27304 = {memory[27304], memory[27305], memory[27306], memory[27307]};
wire [31:0] memory27308 = {memory[27308], memory[27309], memory[27310], memory[27311]};
wire [31:0] memory27312 = {memory[27312], memory[27313], memory[27314], memory[27315]};
wire [31:0] memory27316 = {memory[27316], memory[27317], memory[27318], memory[27319]};
wire [31:0] memory27320 = {memory[27320], memory[27321], memory[27322], memory[27323]};
wire [31:0] memory27324 = {memory[27324], memory[27325], memory[27326], memory[27327]};
wire [31:0] memory27328 = {memory[27328], memory[27329], memory[27330], memory[27331]};
wire [31:0] memory27332 = {memory[27332], memory[27333], memory[27334], memory[27335]};
wire [31:0] memory27336 = {memory[27336], memory[27337], memory[27338], memory[27339]};
wire [31:0] memory27340 = {memory[27340], memory[27341], memory[27342], memory[27343]};
wire [31:0] memory27344 = {memory[27344], memory[27345], memory[27346], memory[27347]};
wire [31:0] memory27348 = {memory[27348], memory[27349], memory[27350], memory[27351]};
wire [31:0] memory27352 = {memory[27352], memory[27353], memory[27354], memory[27355]};
wire [31:0] memory27356 = {memory[27356], memory[27357], memory[27358], memory[27359]};
wire [31:0] memory27360 = {memory[27360], memory[27361], memory[27362], memory[27363]};
wire [31:0] memory27364 = {memory[27364], memory[27365], memory[27366], memory[27367]};
wire [31:0] memory27368 = {memory[27368], memory[27369], memory[27370], memory[27371]};
wire [31:0] memory27372 = {memory[27372], memory[27373], memory[27374], memory[27375]};
wire [31:0] memory27376 = {memory[27376], memory[27377], memory[27378], memory[27379]};
wire [31:0] memory27380 = {memory[27380], memory[27381], memory[27382], memory[27383]};
wire [31:0] memory27384 = {memory[27384], memory[27385], memory[27386], memory[27387]};
wire [31:0] memory27388 = {memory[27388], memory[27389], memory[27390], memory[27391]};
wire [31:0] memory27392 = {memory[27392], memory[27393], memory[27394], memory[27395]};
wire [31:0] memory27396 = {memory[27396], memory[27397], memory[27398], memory[27399]};
wire [31:0] memory27400 = {memory[27400], memory[27401], memory[27402], memory[27403]};
wire [31:0] memory27404 = {memory[27404], memory[27405], memory[27406], memory[27407]};
wire [31:0] memory27408 = {memory[27408], memory[27409], memory[27410], memory[27411]};
wire [31:0] memory27412 = {memory[27412], memory[27413], memory[27414], memory[27415]};
wire [31:0] memory27416 = {memory[27416], memory[27417], memory[27418], memory[27419]};
wire [31:0] memory27420 = {memory[27420], memory[27421], memory[27422], memory[27423]};
wire [31:0] memory27424 = {memory[27424], memory[27425], memory[27426], memory[27427]};
wire [31:0] memory27428 = {memory[27428], memory[27429], memory[27430], memory[27431]};
wire [31:0] memory27432 = {memory[27432], memory[27433], memory[27434], memory[27435]};
wire [31:0] memory27436 = {memory[27436], memory[27437], memory[27438], memory[27439]};
wire [31:0] memory27440 = {memory[27440], memory[27441], memory[27442], memory[27443]};
wire [31:0] memory27444 = {memory[27444], memory[27445], memory[27446], memory[27447]};
wire [31:0] memory27448 = {memory[27448], memory[27449], memory[27450], memory[27451]};
wire [31:0] memory27452 = {memory[27452], memory[27453], memory[27454], memory[27455]};
wire [31:0] memory27456 = {memory[27456], memory[27457], memory[27458], memory[27459]};
wire [31:0] memory27460 = {memory[27460], memory[27461], memory[27462], memory[27463]};
wire [31:0] memory27464 = {memory[27464], memory[27465], memory[27466], memory[27467]};
wire [31:0] memory27468 = {memory[27468], memory[27469], memory[27470], memory[27471]};
wire [31:0] memory27472 = {memory[27472], memory[27473], memory[27474], memory[27475]};
wire [31:0] memory27476 = {memory[27476], memory[27477], memory[27478], memory[27479]};
wire [31:0] memory27480 = {memory[27480], memory[27481], memory[27482], memory[27483]};
wire [31:0] memory27484 = {memory[27484], memory[27485], memory[27486], memory[27487]};
wire [31:0] memory27488 = {memory[27488], memory[27489], memory[27490], memory[27491]};
wire [31:0] memory27492 = {memory[27492], memory[27493], memory[27494], memory[27495]};
wire [31:0] memory27496 = {memory[27496], memory[27497], memory[27498], memory[27499]};
wire [31:0] memory27500 = {memory[27500], memory[27501], memory[27502], memory[27503]};
wire [31:0] memory27504 = {memory[27504], memory[27505], memory[27506], memory[27507]};
wire [31:0] memory27508 = {memory[27508], memory[27509], memory[27510], memory[27511]};
wire [31:0] memory27512 = {memory[27512], memory[27513], memory[27514], memory[27515]};
wire [31:0] memory27516 = {memory[27516], memory[27517], memory[27518], memory[27519]};
wire [31:0] memory27520 = {memory[27520], memory[27521], memory[27522], memory[27523]};
wire [31:0] memory27524 = {memory[27524], memory[27525], memory[27526], memory[27527]};
wire [31:0] memory27528 = {memory[27528], memory[27529], memory[27530], memory[27531]};
wire [31:0] memory27532 = {memory[27532], memory[27533], memory[27534], memory[27535]};
wire [31:0] memory27536 = {memory[27536], memory[27537], memory[27538], memory[27539]};
wire [31:0] memory27540 = {memory[27540], memory[27541], memory[27542], memory[27543]};
wire [31:0] memory27544 = {memory[27544], memory[27545], memory[27546], memory[27547]};
wire [31:0] memory27548 = {memory[27548], memory[27549], memory[27550], memory[27551]};
wire [31:0] memory27552 = {memory[27552], memory[27553], memory[27554], memory[27555]};
wire [31:0] memory27556 = {memory[27556], memory[27557], memory[27558], memory[27559]};
wire [31:0] memory27560 = {memory[27560], memory[27561], memory[27562], memory[27563]};
wire [31:0] memory27564 = {memory[27564], memory[27565], memory[27566], memory[27567]};
wire [31:0] memory27568 = {memory[27568], memory[27569], memory[27570], memory[27571]};
wire [31:0] memory27572 = {memory[27572], memory[27573], memory[27574], memory[27575]};
wire [31:0] memory27576 = {memory[27576], memory[27577], memory[27578], memory[27579]};
wire [31:0] memory27580 = {memory[27580], memory[27581], memory[27582], memory[27583]};
wire [31:0] memory27584 = {memory[27584], memory[27585], memory[27586], memory[27587]};
wire [31:0] memory27588 = {memory[27588], memory[27589], memory[27590], memory[27591]};
wire [31:0] memory27592 = {memory[27592], memory[27593], memory[27594], memory[27595]};
wire [31:0] memory27596 = {memory[27596], memory[27597], memory[27598], memory[27599]};
wire [31:0] memory27600 = {memory[27600], memory[27601], memory[27602], memory[27603]};
wire [31:0] memory27604 = {memory[27604], memory[27605], memory[27606], memory[27607]};
wire [31:0] memory27608 = {memory[27608], memory[27609], memory[27610], memory[27611]};
wire [31:0] memory27612 = {memory[27612], memory[27613], memory[27614], memory[27615]};
wire [31:0] memory27616 = {memory[27616], memory[27617], memory[27618], memory[27619]};
wire [31:0] memory27620 = {memory[27620], memory[27621], memory[27622], memory[27623]};
wire [31:0] memory27624 = {memory[27624], memory[27625], memory[27626], memory[27627]};
wire [31:0] memory27628 = {memory[27628], memory[27629], memory[27630], memory[27631]};
wire [31:0] memory27632 = {memory[27632], memory[27633], memory[27634], memory[27635]};
wire [31:0] memory27636 = {memory[27636], memory[27637], memory[27638], memory[27639]};
wire [31:0] memory27640 = {memory[27640], memory[27641], memory[27642], memory[27643]};
wire [31:0] memory27644 = {memory[27644], memory[27645], memory[27646], memory[27647]};
wire [31:0] memory27648 = {memory[27648], memory[27649], memory[27650], memory[27651]};
wire [31:0] memory27652 = {memory[27652], memory[27653], memory[27654], memory[27655]};
wire [31:0] memory27656 = {memory[27656], memory[27657], memory[27658], memory[27659]};
wire [31:0] memory27660 = {memory[27660], memory[27661], memory[27662], memory[27663]};
wire [31:0] memory27664 = {memory[27664], memory[27665], memory[27666], memory[27667]};
wire [31:0] memory27668 = {memory[27668], memory[27669], memory[27670], memory[27671]};
wire [31:0] memory27672 = {memory[27672], memory[27673], memory[27674], memory[27675]};
wire [31:0] memory27676 = {memory[27676], memory[27677], memory[27678], memory[27679]};
wire [31:0] memory27680 = {memory[27680], memory[27681], memory[27682], memory[27683]};
wire [31:0] memory27684 = {memory[27684], memory[27685], memory[27686], memory[27687]};
wire [31:0] memory27688 = {memory[27688], memory[27689], memory[27690], memory[27691]};
wire [31:0] memory27692 = {memory[27692], memory[27693], memory[27694], memory[27695]};
wire [31:0] memory27696 = {memory[27696], memory[27697], memory[27698], memory[27699]};
wire [31:0] memory27700 = {memory[27700], memory[27701], memory[27702], memory[27703]};
wire [31:0] memory27704 = {memory[27704], memory[27705], memory[27706], memory[27707]};
wire [31:0] memory27708 = {memory[27708], memory[27709], memory[27710], memory[27711]};
wire [31:0] memory27712 = {memory[27712], memory[27713], memory[27714], memory[27715]};
wire [31:0] memory27716 = {memory[27716], memory[27717], memory[27718], memory[27719]};
wire [31:0] memory27720 = {memory[27720], memory[27721], memory[27722], memory[27723]};
wire [31:0] memory27724 = {memory[27724], memory[27725], memory[27726], memory[27727]};
wire [31:0] memory27728 = {memory[27728], memory[27729], memory[27730], memory[27731]};
wire [31:0] memory27732 = {memory[27732], memory[27733], memory[27734], memory[27735]};
wire [31:0] memory27736 = {memory[27736], memory[27737], memory[27738], memory[27739]};
wire [31:0] memory27740 = {memory[27740], memory[27741], memory[27742], memory[27743]};
wire [31:0] memory27744 = {memory[27744], memory[27745], memory[27746], memory[27747]};
wire [31:0] memory27748 = {memory[27748], memory[27749], memory[27750], memory[27751]};
wire [31:0] memory27752 = {memory[27752], memory[27753], memory[27754], memory[27755]};
wire [31:0] memory27756 = {memory[27756], memory[27757], memory[27758], memory[27759]};
wire [31:0] memory27760 = {memory[27760], memory[27761], memory[27762], memory[27763]};
wire [31:0] memory27764 = {memory[27764], memory[27765], memory[27766], memory[27767]};
wire [31:0] memory27768 = {memory[27768], memory[27769], memory[27770], memory[27771]};
wire [31:0] memory27772 = {memory[27772], memory[27773], memory[27774], memory[27775]};
wire [31:0] memory27776 = {memory[27776], memory[27777], memory[27778], memory[27779]};
wire [31:0] memory27780 = {memory[27780], memory[27781], memory[27782], memory[27783]};
wire [31:0] memory27784 = {memory[27784], memory[27785], memory[27786], memory[27787]};
wire [31:0] memory27788 = {memory[27788], memory[27789], memory[27790], memory[27791]};
wire [31:0] memory27792 = {memory[27792], memory[27793], memory[27794], memory[27795]};
wire [31:0] memory27796 = {memory[27796], memory[27797], memory[27798], memory[27799]};
wire [31:0] memory27800 = {memory[27800], memory[27801], memory[27802], memory[27803]};
wire [31:0] memory27804 = {memory[27804], memory[27805], memory[27806], memory[27807]};
wire [31:0] memory27808 = {memory[27808], memory[27809], memory[27810], memory[27811]};
wire [31:0] memory27812 = {memory[27812], memory[27813], memory[27814], memory[27815]};
wire [31:0] memory27816 = {memory[27816], memory[27817], memory[27818], memory[27819]};
wire [31:0] memory27820 = {memory[27820], memory[27821], memory[27822], memory[27823]};
wire [31:0] memory27824 = {memory[27824], memory[27825], memory[27826], memory[27827]};
wire [31:0] memory27828 = {memory[27828], memory[27829], memory[27830], memory[27831]};
wire [31:0] memory27832 = {memory[27832], memory[27833], memory[27834], memory[27835]};
wire [31:0] memory27836 = {memory[27836], memory[27837], memory[27838], memory[27839]};
wire [31:0] memory27840 = {memory[27840], memory[27841], memory[27842], memory[27843]};
wire [31:0] memory27844 = {memory[27844], memory[27845], memory[27846], memory[27847]};
wire [31:0] memory27848 = {memory[27848], memory[27849], memory[27850], memory[27851]};
wire [31:0] memory27852 = {memory[27852], memory[27853], memory[27854], memory[27855]};
wire [31:0] memory27856 = {memory[27856], memory[27857], memory[27858], memory[27859]};
wire [31:0] memory27860 = {memory[27860], memory[27861], memory[27862], memory[27863]};
wire [31:0] memory27864 = {memory[27864], memory[27865], memory[27866], memory[27867]};
wire [31:0] memory27868 = {memory[27868], memory[27869], memory[27870], memory[27871]};
wire [31:0] memory27872 = {memory[27872], memory[27873], memory[27874], memory[27875]};
wire [31:0] memory27876 = {memory[27876], memory[27877], memory[27878], memory[27879]};
wire [31:0] memory27880 = {memory[27880], memory[27881], memory[27882], memory[27883]};
wire [31:0] memory27884 = {memory[27884], memory[27885], memory[27886], memory[27887]};
wire [31:0] memory27888 = {memory[27888], memory[27889], memory[27890], memory[27891]};
wire [31:0] memory27892 = {memory[27892], memory[27893], memory[27894], memory[27895]};
wire [31:0] memory27896 = {memory[27896], memory[27897], memory[27898], memory[27899]};
wire [31:0] memory27900 = {memory[27900], memory[27901], memory[27902], memory[27903]};
wire [31:0] memory27904 = {memory[27904], memory[27905], memory[27906], memory[27907]};
wire [31:0] memory27908 = {memory[27908], memory[27909], memory[27910], memory[27911]};
wire [31:0] memory27912 = {memory[27912], memory[27913], memory[27914], memory[27915]};
wire [31:0] memory27916 = {memory[27916], memory[27917], memory[27918], memory[27919]};
wire [31:0] memory27920 = {memory[27920], memory[27921], memory[27922], memory[27923]};
wire [31:0] memory27924 = {memory[27924], memory[27925], memory[27926], memory[27927]};
wire [31:0] memory27928 = {memory[27928], memory[27929], memory[27930], memory[27931]};
wire [31:0] memory27932 = {memory[27932], memory[27933], memory[27934], memory[27935]};
wire [31:0] memory27936 = {memory[27936], memory[27937], memory[27938], memory[27939]};
wire [31:0] memory27940 = {memory[27940], memory[27941], memory[27942], memory[27943]};
wire [31:0] memory27944 = {memory[27944], memory[27945], memory[27946], memory[27947]};
wire [31:0] memory27948 = {memory[27948], memory[27949], memory[27950], memory[27951]};
wire [31:0] memory27952 = {memory[27952], memory[27953], memory[27954], memory[27955]};
wire [31:0] memory27956 = {memory[27956], memory[27957], memory[27958], memory[27959]};
wire [31:0] memory27960 = {memory[27960], memory[27961], memory[27962], memory[27963]};
wire [31:0] memory27964 = {memory[27964], memory[27965], memory[27966], memory[27967]};
wire [31:0] memory27968 = {memory[27968], memory[27969], memory[27970], memory[27971]};
wire [31:0] memory27972 = {memory[27972], memory[27973], memory[27974], memory[27975]};
wire [31:0] memory27976 = {memory[27976], memory[27977], memory[27978], memory[27979]};
wire [31:0] memory27980 = {memory[27980], memory[27981], memory[27982], memory[27983]};
wire [31:0] memory27984 = {memory[27984], memory[27985], memory[27986], memory[27987]};
wire [31:0] memory27988 = {memory[27988], memory[27989], memory[27990], memory[27991]};
wire [31:0] memory27992 = {memory[27992], memory[27993], memory[27994], memory[27995]};
wire [31:0] memory27996 = {memory[27996], memory[27997], memory[27998], memory[27999]};
wire [31:0] memory28000 = {memory[28000], memory[28001], memory[28002], memory[28003]};
wire [31:0] memory28004 = {memory[28004], memory[28005], memory[28006], memory[28007]};
wire [31:0] memory28008 = {memory[28008], memory[28009], memory[28010], memory[28011]};
wire [31:0] memory28012 = {memory[28012], memory[28013], memory[28014], memory[28015]};
wire [31:0] memory28016 = {memory[28016], memory[28017], memory[28018], memory[28019]};
wire [31:0] memory28020 = {memory[28020], memory[28021], memory[28022], memory[28023]};
wire [31:0] memory28024 = {memory[28024], memory[28025], memory[28026], memory[28027]};
wire [31:0] memory28028 = {memory[28028], memory[28029], memory[28030], memory[28031]};
wire [31:0] memory28032 = {memory[28032], memory[28033], memory[28034], memory[28035]};
wire [31:0] memory28036 = {memory[28036], memory[28037], memory[28038], memory[28039]};
wire [31:0] memory28040 = {memory[28040], memory[28041], memory[28042], memory[28043]};
wire [31:0] memory28044 = {memory[28044], memory[28045], memory[28046], memory[28047]};
wire [31:0] memory28048 = {memory[28048], memory[28049], memory[28050], memory[28051]};
wire [31:0] memory28052 = {memory[28052], memory[28053], memory[28054], memory[28055]};
wire [31:0] memory28056 = {memory[28056], memory[28057], memory[28058], memory[28059]};
wire [31:0] memory28060 = {memory[28060], memory[28061], memory[28062], memory[28063]};
wire [31:0] memory28064 = {memory[28064], memory[28065], memory[28066], memory[28067]};
wire [31:0] memory28068 = {memory[28068], memory[28069], memory[28070], memory[28071]};
wire [31:0] memory28072 = {memory[28072], memory[28073], memory[28074], memory[28075]};
wire [31:0] memory28076 = {memory[28076], memory[28077], memory[28078], memory[28079]};
wire [31:0] memory28080 = {memory[28080], memory[28081], memory[28082], memory[28083]};
wire [31:0] memory28084 = {memory[28084], memory[28085], memory[28086], memory[28087]};
wire [31:0] memory28088 = {memory[28088], memory[28089], memory[28090], memory[28091]};
wire [31:0] memory28092 = {memory[28092], memory[28093], memory[28094], memory[28095]};
wire [31:0] memory28096 = {memory[28096], memory[28097], memory[28098], memory[28099]};
wire [31:0] memory28100 = {memory[28100], memory[28101], memory[28102], memory[28103]};
wire [31:0] memory28104 = {memory[28104], memory[28105], memory[28106], memory[28107]};
wire [31:0] memory28108 = {memory[28108], memory[28109], memory[28110], memory[28111]};
wire [31:0] memory28112 = {memory[28112], memory[28113], memory[28114], memory[28115]};
wire [31:0] memory28116 = {memory[28116], memory[28117], memory[28118], memory[28119]};
wire [31:0] memory28120 = {memory[28120], memory[28121], memory[28122], memory[28123]};
wire [31:0] memory28124 = {memory[28124], memory[28125], memory[28126], memory[28127]};
wire [31:0] memory28128 = {memory[28128], memory[28129], memory[28130], memory[28131]};
wire [31:0] memory28132 = {memory[28132], memory[28133], memory[28134], memory[28135]};
wire [31:0] memory28136 = {memory[28136], memory[28137], memory[28138], memory[28139]};
wire [31:0] memory28140 = {memory[28140], memory[28141], memory[28142], memory[28143]};
wire [31:0] memory28144 = {memory[28144], memory[28145], memory[28146], memory[28147]};
wire [31:0] memory28148 = {memory[28148], memory[28149], memory[28150], memory[28151]};
wire [31:0] memory28152 = {memory[28152], memory[28153], memory[28154], memory[28155]};
wire [31:0] memory28156 = {memory[28156], memory[28157], memory[28158], memory[28159]};
wire [31:0] memory28160 = {memory[28160], memory[28161], memory[28162], memory[28163]};
wire [31:0] memory28164 = {memory[28164], memory[28165], memory[28166], memory[28167]};
wire [31:0] memory28168 = {memory[28168], memory[28169], memory[28170], memory[28171]};
wire [31:0] memory28172 = {memory[28172], memory[28173], memory[28174], memory[28175]};
wire [31:0] memory28176 = {memory[28176], memory[28177], memory[28178], memory[28179]};
wire [31:0] memory28180 = {memory[28180], memory[28181], memory[28182], memory[28183]};
wire [31:0] memory28184 = {memory[28184], memory[28185], memory[28186], memory[28187]};
wire [31:0] memory28188 = {memory[28188], memory[28189], memory[28190], memory[28191]};
wire [31:0] memory28192 = {memory[28192], memory[28193], memory[28194], memory[28195]};
wire [31:0] memory28196 = {memory[28196], memory[28197], memory[28198], memory[28199]};
wire [31:0] memory28200 = {memory[28200], memory[28201], memory[28202], memory[28203]};
wire [31:0] memory28204 = {memory[28204], memory[28205], memory[28206], memory[28207]};
wire [31:0] memory28208 = {memory[28208], memory[28209], memory[28210], memory[28211]};
wire [31:0] memory28212 = {memory[28212], memory[28213], memory[28214], memory[28215]};
wire [31:0] memory28216 = {memory[28216], memory[28217], memory[28218], memory[28219]};
wire [31:0] memory28220 = {memory[28220], memory[28221], memory[28222], memory[28223]};
wire [31:0] memory28224 = {memory[28224], memory[28225], memory[28226], memory[28227]};
wire [31:0] memory28228 = {memory[28228], memory[28229], memory[28230], memory[28231]};
wire [31:0] memory28232 = {memory[28232], memory[28233], memory[28234], memory[28235]};
wire [31:0] memory28236 = {memory[28236], memory[28237], memory[28238], memory[28239]};
wire [31:0] memory28240 = {memory[28240], memory[28241], memory[28242], memory[28243]};
wire [31:0] memory28244 = {memory[28244], memory[28245], memory[28246], memory[28247]};
wire [31:0] memory28248 = {memory[28248], memory[28249], memory[28250], memory[28251]};
wire [31:0] memory28252 = {memory[28252], memory[28253], memory[28254], memory[28255]};
wire [31:0] memory28256 = {memory[28256], memory[28257], memory[28258], memory[28259]};
wire [31:0] memory28260 = {memory[28260], memory[28261], memory[28262], memory[28263]};
wire [31:0] memory28264 = {memory[28264], memory[28265], memory[28266], memory[28267]};
wire [31:0] memory28268 = {memory[28268], memory[28269], memory[28270], memory[28271]};
wire [31:0] memory28272 = {memory[28272], memory[28273], memory[28274], memory[28275]};
wire [31:0] memory28276 = {memory[28276], memory[28277], memory[28278], memory[28279]};
wire [31:0] memory28280 = {memory[28280], memory[28281], memory[28282], memory[28283]};
wire [31:0] memory28284 = {memory[28284], memory[28285], memory[28286], memory[28287]};
wire [31:0] memory28288 = {memory[28288], memory[28289], memory[28290], memory[28291]};
wire [31:0] memory28292 = {memory[28292], memory[28293], memory[28294], memory[28295]};
wire [31:0] memory28296 = {memory[28296], memory[28297], memory[28298], memory[28299]};
wire [31:0] memory28300 = {memory[28300], memory[28301], memory[28302], memory[28303]};
wire [31:0] memory28304 = {memory[28304], memory[28305], memory[28306], memory[28307]};
wire [31:0] memory28308 = {memory[28308], memory[28309], memory[28310], memory[28311]};
wire [31:0] memory28312 = {memory[28312], memory[28313], memory[28314], memory[28315]};
wire [31:0] memory28316 = {memory[28316], memory[28317], memory[28318], memory[28319]};
wire [31:0] memory28320 = {memory[28320], memory[28321], memory[28322], memory[28323]};
wire [31:0] memory28324 = {memory[28324], memory[28325], memory[28326], memory[28327]};
wire [31:0] memory28328 = {memory[28328], memory[28329], memory[28330], memory[28331]};
wire [31:0] memory28332 = {memory[28332], memory[28333], memory[28334], memory[28335]};
wire [31:0] memory28336 = {memory[28336], memory[28337], memory[28338], memory[28339]};
wire [31:0] memory28340 = {memory[28340], memory[28341], memory[28342], memory[28343]};
wire [31:0] memory28344 = {memory[28344], memory[28345], memory[28346], memory[28347]};
wire [31:0] memory28348 = {memory[28348], memory[28349], memory[28350], memory[28351]};
wire [31:0] memory28352 = {memory[28352], memory[28353], memory[28354], memory[28355]};
wire [31:0] memory28356 = {memory[28356], memory[28357], memory[28358], memory[28359]};
wire [31:0] memory28360 = {memory[28360], memory[28361], memory[28362], memory[28363]};
wire [31:0] memory28364 = {memory[28364], memory[28365], memory[28366], memory[28367]};
wire [31:0] memory28368 = {memory[28368], memory[28369], memory[28370], memory[28371]};
wire [31:0] memory28372 = {memory[28372], memory[28373], memory[28374], memory[28375]};
wire [31:0] memory28376 = {memory[28376], memory[28377], memory[28378], memory[28379]};
wire [31:0] memory28380 = {memory[28380], memory[28381], memory[28382], memory[28383]};
wire [31:0] memory28384 = {memory[28384], memory[28385], memory[28386], memory[28387]};
wire [31:0] memory28388 = {memory[28388], memory[28389], memory[28390], memory[28391]};
wire [31:0] memory28392 = {memory[28392], memory[28393], memory[28394], memory[28395]};
wire [31:0] memory28396 = {memory[28396], memory[28397], memory[28398], memory[28399]};
wire [31:0] memory28400 = {memory[28400], memory[28401], memory[28402], memory[28403]};
wire [31:0] memory28404 = {memory[28404], memory[28405], memory[28406], memory[28407]};
wire [31:0] memory28408 = {memory[28408], memory[28409], memory[28410], memory[28411]};
wire [31:0] memory28412 = {memory[28412], memory[28413], memory[28414], memory[28415]};
wire [31:0] memory28416 = {memory[28416], memory[28417], memory[28418], memory[28419]};
wire [31:0] memory28420 = {memory[28420], memory[28421], memory[28422], memory[28423]};
wire [31:0] memory28424 = {memory[28424], memory[28425], memory[28426], memory[28427]};
wire [31:0] memory28428 = {memory[28428], memory[28429], memory[28430], memory[28431]};
wire [31:0] memory28432 = {memory[28432], memory[28433], memory[28434], memory[28435]};
wire [31:0] memory28436 = {memory[28436], memory[28437], memory[28438], memory[28439]};
wire [31:0] memory28440 = {memory[28440], memory[28441], memory[28442], memory[28443]};
wire [31:0] memory28444 = {memory[28444], memory[28445], memory[28446], memory[28447]};
wire [31:0] memory28448 = {memory[28448], memory[28449], memory[28450], memory[28451]};
wire [31:0] memory28452 = {memory[28452], memory[28453], memory[28454], memory[28455]};
wire [31:0] memory28456 = {memory[28456], memory[28457], memory[28458], memory[28459]};
wire [31:0] memory28460 = {memory[28460], memory[28461], memory[28462], memory[28463]};
wire [31:0] memory28464 = {memory[28464], memory[28465], memory[28466], memory[28467]};
wire [31:0] memory28468 = {memory[28468], memory[28469], memory[28470], memory[28471]};
wire [31:0] memory28472 = {memory[28472], memory[28473], memory[28474], memory[28475]};
wire [31:0] memory28476 = {memory[28476], memory[28477], memory[28478], memory[28479]};
wire [31:0] memory28480 = {memory[28480], memory[28481], memory[28482], memory[28483]};
wire [31:0] memory28484 = {memory[28484], memory[28485], memory[28486], memory[28487]};
wire [31:0] memory28488 = {memory[28488], memory[28489], memory[28490], memory[28491]};
wire [31:0] memory28492 = {memory[28492], memory[28493], memory[28494], memory[28495]};
wire [31:0] memory28496 = {memory[28496], memory[28497], memory[28498], memory[28499]};
wire [31:0] memory28500 = {memory[28500], memory[28501], memory[28502], memory[28503]};
wire [31:0] memory28504 = {memory[28504], memory[28505], memory[28506], memory[28507]};
wire [31:0] memory28508 = {memory[28508], memory[28509], memory[28510], memory[28511]};
wire [31:0] memory28512 = {memory[28512], memory[28513], memory[28514], memory[28515]};
wire [31:0] memory28516 = {memory[28516], memory[28517], memory[28518], memory[28519]};
wire [31:0] memory28520 = {memory[28520], memory[28521], memory[28522], memory[28523]};
wire [31:0] memory28524 = {memory[28524], memory[28525], memory[28526], memory[28527]};
wire [31:0] memory28528 = {memory[28528], memory[28529], memory[28530], memory[28531]};
wire [31:0] memory28532 = {memory[28532], memory[28533], memory[28534], memory[28535]};
wire [31:0] memory28536 = {memory[28536], memory[28537], memory[28538], memory[28539]};
wire [31:0] memory28540 = {memory[28540], memory[28541], memory[28542], memory[28543]};
wire [31:0] memory28544 = {memory[28544], memory[28545], memory[28546], memory[28547]};
wire [31:0] memory28548 = {memory[28548], memory[28549], memory[28550], memory[28551]};
wire [31:0] memory28552 = {memory[28552], memory[28553], memory[28554], memory[28555]};
wire [31:0] memory28556 = {memory[28556], memory[28557], memory[28558], memory[28559]};
wire [31:0] memory28560 = {memory[28560], memory[28561], memory[28562], memory[28563]};
wire [31:0] memory28564 = {memory[28564], memory[28565], memory[28566], memory[28567]};
wire [31:0] memory28568 = {memory[28568], memory[28569], memory[28570], memory[28571]};
wire [31:0] memory28572 = {memory[28572], memory[28573], memory[28574], memory[28575]};
wire [31:0] memory28576 = {memory[28576], memory[28577], memory[28578], memory[28579]};
wire [31:0] memory28580 = {memory[28580], memory[28581], memory[28582], memory[28583]};
wire [31:0] memory28584 = {memory[28584], memory[28585], memory[28586], memory[28587]};
wire [31:0] memory28588 = {memory[28588], memory[28589], memory[28590], memory[28591]};
wire [31:0] memory28592 = {memory[28592], memory[28593], memory[28594], memory[28595]};
wire [31:0] memory28596 = {memory[28596], memory[28597], memory[28598], memory[28599]};
wire [31:0] memory28600 = {memory[28600], memory[28601], memory[28602], memory[28603]};
wire [31:0] memory28604 = {memory[28604], memory[28605], memory[28606], memory[28607]};
wire [31:0] memory28608 = {memory[28608], memory[28609], memory[28610], memory[28611]};
wire [31:0] memory28612 = {memory[28612], memory[28613], memory[28614], memory[28615]};
wire [31:0] memory28616 = {memory[28616], memory[28617], memory[28618], memory[28619]};
wire [31:0] memory28620 = {memory[28620], memory[28621], memory[28622], memory[28623]};
wire [31:0] memory28624 = {memory[28624], memory[28625], memory[28626], memory[28627]};
wire [31:0] memory28628 = {memory[28628], memory[28629], memory[28630], memory[28631]};
wire [31:0] memory28632 = {memory[28632], memory[28633], memory[28634], memory[28635]};
wire [31:0] memory28636 = {memory[28636], memory[28637], memory[28638], memory[28639]};
wire [31:0] memory28640 = {memory[28640], memory[28641], memory[28642], memory[28643]};
wire [31:0] memory28644 = {memory[28644], memory[28645], memory[28646], memory[28647]};
wire [31:0] memory28648 = {memory[28648], memory[28649], memory[28650], memory[28651]};
wire [31:0] memory28652 = {memory[28652], memory[28653], memory[28654], memory[28655]};
wire [31:0] memory28656 = {memory[28656], memory[28657], memory[28658], memory[28659]};
wire [31:0] memory28660 = {memory[28660], memory[28661], memory[28662], memory[28663]};
wire [31:0] memory28664 = {memory[28664], memory[28665], memory[28666], memory[28667]};
wire [31:0] memory28668 = {memory[28668], memory[28669], memory[28670], memory[28671]};
wire [31:0] memory28672 = {memory[28672], memory[28673], memory[28674], memory[28675]};
wire [31:0] memory28676 = {memory[28676], memory[28677], memory[28678], memory[28679]};
wire [31:0] memory28680 = {memory[28680], memory[28681], memory[28682], memory[28683]};
wire [31:0] memory28684 = {memory[28684], memory[28685], memory[28686], memory[28687]};
wire [31:0] memory28688 = {memory[28688], memory[28689], memory[28690], memory[28691]};
wire [31:0] memory28692 = {memory[28692], memory[28693], memory[28694], memory[28695]};
wire [31:0] memory28696 = {memory[28696], memory[28697], memory[28698], memory[28699]};
wire [31:0] memory28700 = {memory[28700], memory[28701], memory[28702], memory[28703]};
wire [31:0] memory28704 = {memory[28704], memory[28705], memory[28706], memory[28707]};
wire [31:0] memory28708 = {memory[28708], memory[28709], memory[28710], memory[28711]};
wire [31:0] memory28712 = {memory[28712], memory[28713], memory[28714], memory[28715]};
wire [31:0] memory28716 = {memory[28716], memory[28717], memory[28718], memory[28719]};
wire [31:0] memory28720 = {memory[28720], memory[28721], memory[28722], memory[28723]};
wire [31:0] memory28724 = {memory[28724], memory[28725], memory[28726], memory[28727]};
wire [31:0] memory28728 = {memory[28728], memory[28729], memory[28730], memory[28731]};
wire [31:0] memory28732 = {memory[28732], memory[28733], memory[28734], memory[28735]};
wire [31:0] memory28736 = {memory[28736], memory[28737], memory[28738], memory[28739]};
wire [31:0] memory28740 = {memory[28740], memory[28741], memory[28742], memory[28743]};
wire [31:0] memory28744 = {memory[28744], memory[28745], memory[28746], memory[28747]};
wire [31:0] memory28748 = {memory[28748], memory[28749], memory[28750], memory[28751]};
wire [31:0] memory28752 = {memory[28752], memory[28753], memory[28754], memory[28755]};
wire [31:0] memory28756 = {memory[28756], memory[28757], memory[28758], memory[28759]};
wire [31:0] memory28760 = {memory[28760], memory[28761], memory[28762], memory[28763]};
wire [31:0] memory28764 = {memory[28764], memory[28765], memory[28766], memory[28767]};
wire [31:0] memory28768 = {memory[28768], memory[28769], memory[28770], memory[28771]};
wire [31:0] memory28772 = {memory[28772], memory[28773], memory[28774], memory[28775]};
wire [31:0] memory28776 = {memory[28776], memory[28777], memory[28778], memory[28779]};
wire [31:0] memory28780 = {memory[28780], memory[28781], memory[28782], memory[28783]};
wire [31:0] memory28784 = {memory[28784], memory[28785], memory[28786], memory[28787]};
wire [31:0] memory28788 = {memory[28788], memory[28789], memory[28790], memory[28791]};
wire [31:0] memory28792 = {memory[28792], memory[28793], memory[28794], memory[28795]};
wire [31:0] memory28796 = {memory[28796], memory[28797], memory[28798], memory[28799]};
wire [31:0] memory28800 = {memory[28800], memory[28801], memory[28802], memory[28803]};
wire [31:0] memory28804 = {memory[28804], memory[28805], memory[28806], memory[28807]};
wire [31:0] memory28808 = {memory[28808], memory[28809], memory[28810], memory[28811]};
wire [31:0] memory28812 = {memory[28812], memory[28813], memory[28814], memory[28815]};
wire [31:0] memory28816 = {memory[28816], memory[28817], memory[28818], memory[28819]};
wire [31:0] memory28820 = {memory[28820], memory[28821], memory[28822], memory[28823]};
wire [31:0] memory28824 = {memory[28824], memory[28825], memory[28826], memory[28827]};
wire [31:0] memory28828 = {memory[28828], memory[28829], memory[28830], memory[28831]};
wire [31:0] memory28832 = {memory[28832], memory[28833], memory[28834], memory[28835]};
wire [31:0] memory28836 = {memory[28836], memory[28837], memory[28838], memory[28839]};
wire [31:0] memory28840 = {memory[28840], memory[28841], memory[28842], memory[28843]};
wire [31:0] memory28844 = {memory[28844], memory[28845], memory[28846], memory[28847]};
wire [31:0] memory28848 = {memory[28848], memory[28849], memory[28850], memory[28851]};
wire [31:0] memory28852 = {memory[28852], memory[28853], memory[28854], memory[28855]};
wire [31:0] memory28856 = {memory[28856], memory[28857], memory[28858], memory[28859]};
wire [31:0] memory28860 = {memory[28860], memory[28861], memory[28862], memory[28863]};
wire [31:0] memory28864 = {memory[28864], memory[28865], memory[28866], memory[28867]};
wire [31:0] memory28868 = {memory[28868], memory[28869], memory[28870], memory[28871]};
wire [31:0] memory28872 = {memory[28872], memory[28873], memory[28874], memory[28875]};
wire [31:0] memory28876 = {memory[28876], memory[28877], memory[28878], memory[28879]};
wire [31:0] memory28880 = {memory[28880], memory[28881], memory[28882], memory[28883]};
wire [31:0] memory28884 = {memory[28884], memory[28885], memory[28886], memory[28887]};
wire [31:0] memory28888 = {memory[28888], memory[28889], memory[28890], memory[28891]};
wire [31:0] memory28892 = {memory[28892], memory[28893], memory[28894], memory[28895]};
wire [31:0] memory28896 = {memory[28896], memory[28897], memory[28898], memory[28899]};
wire [31:0] memory28900 = {memory[28900], memory[28901], memory[28902], memory[28903]};
wire [31:0] memory28904 = {memory[28904], memory[28905], memory[28906], memory[28907]};
wire [31:0] memory28908 = {memory[28908], memory[28909], memory[28910], memory[28911]};
wire [31:0] memory28912 = {memory[28912], memory[28913], memory[28914], memory[28915]};
wire [31:0] memory28916 = {memory[28916], memory[28917], memory[28918], memory[28919]};
wire [31:0] memory28920 = {memory[28920], memory[28921], memory[28922], memory[28923]};
wire [31:0] memory28924 = {memory[28924], memory[28925], memory[28926], memory[28927]};
wire [31:0] memory28928 = {memory[28928], memory[28929], memory[28930], memory[28931]};
wire [31:0] memory28932 = {memory[28932], memory[28933], memory[28934], memory[28935]};
wire [31:0] memory28936 = {memory[28936], memory[28937], memory[28938], memory[28939]};
wire [31:0] memory28940 = {memory[28940], memory[28941], memory[28942], memory[28943]};
wire [31:0] memory28944 = {memory[28944], memory[28945], memory[28946], memory[28947]};
wire [31:0] memory28948 = {memory[28948], memory[28949], memory[28950], memory[28951]};
wire [31:0] memory28952 = {memory[28952], memory[28953], memory[28954], memory[28955]};
wire [31:0] memory28956 = {memory[28956], memory[28957], memory[28958], memory[28959]};
wire [31:0] memory28960 = {memory[28960], memory[28961], memory[28962], memory[28963]};
wire [31:0] memory28964 = {memory[28964], memory[28965], memory[28966], memory[28967]};
wire [31:0] memory28968 = {memory[28968], memory[28969], memory[28970], memory[28971]};
wire [31:0] memory28972 = {memory[28972], memory[28973], memory[28974], memory[28975]};
wire [31:0] memory28976 = {memory[28976], memory[28977], memory[28978], memory[28979]};
wire [31:0] memory28980 = {memory[28980], memory[28981], memory[28982], memory[28983]};
wire [31:0] memory28984 = {memory[28984], memory[28985], memory[28986], memory[28987]};
wire [31:0] memory28988 = {memory[28988], memory[28989], memory[28990], memory[28991]};
wire [31:0] memory28992 = {memory[28992], memory[28993], memory[28994], memory[28995]};
wire [31:0] memory28996 = {memory[28996], memory[28997], memory[28998], memory[28999]};
wire [31:0] memory29000 = {memory[29000], memory[29001], memory[29002], memory[29003]};
wire [31:0] memory29004 = {memory[29004], memory[29005], memory[29006], memory[29007]};
wire [31:0] memory29008 = {memory[29008], memory[29009], memory[29010], memory[29011]};
wire [31:0] memory29012 = {memory[29012], memory[29013], memory[29014], memory[29015]};
wire [31:0] memory29016 = {memory[29016], memory[29017], memory[29018], memory[29019]};
wire [31:0] memory29020 = {memory[29020], memory[29021], memory[29022], memory[29023]};
wire [31:0] memory29024 = {memory[29024], memory[29025], memory[29026], memory[29027]};
wire [31:0] memory29028 = {memory[29028], memory[29029], memory[29030], memory[29031]};
wire [31:0] memory29032 = {memory[29032], memory[29033], memory[29034], memory[29035]};
wire [31:0] memory29036 = {memory[29036], memory[29037], memory[29038], memory[29039]};
wire [31:0] memory29040 = {memory[29040], memory[29041], memory[29042], memory[29043]};
wire [31:0] memory29044 = {memory[29044], memory[29045], memory[29046], memory[29047]};
wire [31:0] memory29048 = {memory[29048], memory[29049], memory[29050], memory[29051]};
wire [31:0] memory29052 = {memory[29052], memory[29053], memory[29054], memory[29055]};
wire [31:0] memory29056 = {memory[29056], memory[29057], memory[29058], memory[29059]};
wire [31:0] memory29060 = {memory[29060], memory[29061], memory[29062], memory[29063]};
wire [31:0] memory29064 = {memory[29064], memory[29065], memory[29066], memory[29067]};
wire [31:0] memory29068 = {memory[29068], memory[29069], memory[29070], memory[29071]};
wire [31:0] memory29072 = {memory[29072], memory[29073], memory[29074], memory[29075]};
wire [31:0] memory29076 = {memory[29076], memory[29077], memory[29078], memory[29079]};
wire [31:0] memory29080 = {memory[29080], memory[29081], memory[29082], memory[29083]};
wire [31:0] memory29084 = {memory[29084], memory[29085], memory[29086], memory[29087]};
wire [31:0] memory29088 = {memory[29088], memory[29089], memory[29090], memory[29091]};
wire [31:0] memory29092 = {memory[29092], memory[29093], memory[29094], memory[29095]};
wire [31:0] memory29096 = {memory[29096], memory[29097], memory[29098], memory[29099]};
wire [31:0] memory29100 = {memory[29100], memory[29101], memory[29102], memory[29103]};
wire [31:0] memory29104 = {memory[29104], memory[29105], memory[29106], memory[29107]};
wire [31:0] memory29108 = {memory[29108], memory[29109], memory[29110], memory[29111]};
wire [31:0] memory29112 = {memory[29112], memory[29113], memory[29114], memory[29115]};
wire [31:0] memory29116 = {memory[29116], memory[29117], memory[29118], memory[29119]};
wire [31:0] memory29120 = {memory[29120], memory[29121], memory[29122], memory[29123]};
wire [31:0] memory29124 = {memory[29124], memory[29125], memory[29126], memory[29127]};
wire [31:0] memory29128 = {memory[29128], memory[29129], memory[29130], memory[29131]};
wire [31:0] memory29132 = {memory[29132], memory[29133], memory[29134], memory[29135]};
wire [31:0] memory29136 = {memory[29136], memory[29137], memory[29138], memory[29139]};
wire [31:0] memory29140 = {memory[29140], memory[29141], memory[29142], memory[29143]};
wire [31:0] memory29144 = {memory[29144], memory[29145], memory[29146], memory[29147]};
wire [31:0] memory29148 = {memory[29148], memory[29149], memory[29150], memory[29151]};
wire [31:0] memory29152 = {memory[29152], memory[29153], memory[29154], memory[29155]};
wire [31:0] memory29156 = {memory[29156], memory[29157], memory[29158], memory[29159]};
wire [31:0] memory29160 = {memory[29160], memory[29161], memory[29162], memory[29163]};
wire [31:0] memory29164 = {memory[29164], memory[29165], memory[29166], memory[29167]};
wire [31:0] memory29168 = {memory[29168], memory[29169], memory[29170], memory[29171]};
wire [31:0] memory29172 = {memory[29172], memory[29173], memory[29174], memory[29175]};
wire [31:0] memory29176 = {memory[29176], memory[29177], memory[29178], memory[29179]};
wire [31:0] memory29180 = {memory[29180], memory[29181], memory[29182], memory[29183]};
wire [31:0] memory29184 = {memory[29184], memory[29185], memory[29186], memory[29187]};
wire [31:0] memory29188 = {memory[29188], memory[29189], memory[29190], memory[29191]};
wire [31:0] memory29192 = {memory[29192], memory[29193], memory[29194], memory[29195]};
wire [31:0] memory29196 = {memory[29196], memory[29197], memory[29198], memory[29199]};
wire [31:0] memory29200 = {memory[29200], memory[29201], memory[29202], memory[29203]};
wire [31:0] memory29204 = {memory[29204], memory[29205], memory[29206], memory[29207]};
wire [31:0] memory29208 = {memory[29208], memory[29209], memory[29210], memory[29211]};
wire [31:0] memory29212 = {memory[29212], memory[29213], memory[29214], memory[29215]};
wire [31:0] memory29216 = {memory[29216], memory[29217], memory[29218], memory[29219]};
wire [31:0] memory29220 = {memory[29220], memory[29221], memory[29222], memory[29223]};
wire [31:0] memory29224 = {memory[29224], memory[29225], memory[29226], memory[29227]};
wire [31:0] memory29228 = {memory[29228], memory[29229], memory[29230], memory[29231]};
wire [31:0] memory29232 = {memory[29232], memory[29233], memory[29234], memory[29235]};
wire [31:0] memory29236 = {memory[29236], memory[29237], memory[29238], memory[29239]};
wire [31:0] memory29240 = {memory[29240], memory[29241], memory[29242], memory[29243]};
wire [31:0] memory29244 = {memory[29244], memory[29245], memory[29246], memory[29247]};
wire [31:0] memory29248 = {memory[29248], memory[29249], memory[29250], memory[29251]};
wire [31:0] memory29252 = {memory[29252], memory[29253], memory[29254], memory[29255]};
wire [31:0] memory29256 = {memory[29256], memory[29257], memory[29258], memory[29259]};
wire [31:0] memory29260 = {memory[29260], memory[29261], memory[29262], memory[29263]};
wire [31:0] memory29264 = {memory[29264], memory[29265], memory[29266], memory[29267]};
wire [31:0] memory29268 = {memory[29268], memory[29269], memory[29270], memory[29271]};
wire [31:0] memory29272 = {memory[29272], memory[29273], memory[29274], memory[29275]};
wire [31:0] memory29276 = {memory[29276], memory[29277], memory[29278], memory[29279]};
wire [31:0] memory29280 = {memory[29280], memory[29281], memory[29282], memory[29283]};
wire [31:0] memory29284 = {memory[29284], memory[29285], memory[29286], memory[29287]};
wire [31:0] memory29288 = {memory[29288], memory[29289], memory[29290], memory[29291]};
wire [31:0] memory29292 = {memory[29292], memory[29293], memory[29294], memory[29295]};
wire [31:0] memory29296 = {memory[29296], memory[29297], memory[29298], memory[29299]};
wire [31:0] memory29300 = {memory[29300], memory[29301], memory[29302], memory[29303]};
wire [31:0] memory29304 = {memory[29304], memory[29305], memory[29306], memory[29307]};
wire [31:0] memory29308 = {memory[29308], memory[29309], memory[29310], memory[29311]};
wire [31:0] memory29312 = {memory[29312], memory[29313], memory[29314], memory[29315]};
wire [31:0] memory29316 = {memory[29316], memory[29317], memory[29318], memory[29319]};
wire [31:0] memory29320 = {memory[29320], memory[29321], memory[29322], memory[29323]};
wire [31:0] memory29324 = {memory[29324], memory[29325], memory[29326], memory[29327]};
wire [31:0] memory29328 = {memory[29328], memory[29329], memory[29330], memory[29331]};
wire [31:0] memory29332 = {memory[29332], memory[29333], memory[29334], memory[29335]};
wire [31:0] memory29336 = {memory[29336], memory[29337], memory[29338], memory[29339]};
wire [31:0] memory29340 = {memory[29340], memory[29341], memory[29342], memory[29343]};
wire [31:0] memory29344 = {memory[29344], memory[29345], memory[29346], memory[29347]};
wire [31:0] memory29348 = {memory[29348], memory[29349], memory[29350], memory[29351]};
wire [31:0] memory29352 = {memory[29352], memory[29353], memory[29354], memory[29355]};
wire [31:0] memory29356 = {memory[29356], memory[29357], memory[29358], memory[29359]};
wire [31:0] memory29360 = {memory[29360], memory[29361], memory[29362], memory[29363]};
wire [31:0] memory29364 = {memory[29364], memory[29365], memory[29366], memory[29367]};
wire [31:0] memory29368 = {memory[29368], memory[29369], memory[29370], memory[29371]};
wire [31:0] memory29372 = {memory[29372], memory[29373], memory[29374], memory[29375]};
wire [31:0] memory29376 = {memory[29376], memory[29377], memory[29378], memory[29379]};
wire [31:0] memory29380 = {memory[29380], memory[29381], memory[29382], memory[29383]};
wire [31:0] memory29384 = {memory[29384], memory[29385], memory[29386], memory[29387]};
wire [31:0] memory29388 = {memory[29388], memory[29389], memory[29390], memory[29391]};
wire [31:0] memory29392 = {memory[29392], memory[29393], memory[29394], memory[29395]};
wire [31:0] memory29396 = {memory[29396], memory[29397], memory[29398], memory[29399]};
wire [31:0] memory29400 = {memory[29400], memory[29401], memory[29402], memory[29403]};
wire [31:0] memory29404 = {memory[29404], memory[29405], memory[29406], memory[29407]};
wire [31:0] memory29408 = {memory[29408], memory[29409], memory[29410], memory[29411]};
wire [31:0] memory29412 = {memory[29412], memory[29413], memory[29414], memory[29415]};
wire [31:0] memory29416 = {memory[29416], memory[29417], memory[29418], memory[29419]};
wire [31:0] memory29420 = {memory[29420], memory[29421], memory[29422], memory[29423]};
wire [31:0] memory29424 = {memory[29424], memory[29425], memory[29426], memory[29427]};
wire [31:0] memory29428 = {memory[29428], memory[29429], memory[29430], memory[29431]};
wire [31:0] memory29432 = {memory[29432], memory[29433], memory[29434], memory[29435]};
wire [31:0] memory29436 = {memory[29436], memory[29437], memory[29438], memory[29439]};
wire [31:0] memory29440 = {memory[29440], memory[29441], memory[29442], memory[29443]};
wire [31:0] memory29444 = {memory[29444], memory[29445], memory[29446], memory[29447]};
wire [31:0] memory29448 = {memory[29448], memory[29449], memory[29450], memory[29451]};
wire [31:0] memory29452 = {memory[29452], memory[29453], memory[29454], memory[29455]};
wire [31:0] memory29456 = {memory[29456], memory[29457], memory[29458], memory[29459]};
wire [31:0] memory29460 = {memory[29460], memory[29461], memory[29462], memory[29463]};
wire [31:0] memory29464 = {memory[29464], memory[29465], memory[29466], memory[29467]};
wire [31:0] memory29468 = {memory[29468], memory[29469], memory[29470], memory[29471]};
wire [31:0] memory29472 = {memory[29472], memory[29473], memory[29474], memory[29475]};
wire [31:0] memory29476 = {memory[29476], memory[29477], memory[29478], memory[29479]};
wire [31:0] memory29480 = {memory[29480], memory[29481], memory[29482], memory[29483]};
wire [31:0] memory29484 = {memory[29484], memory[29485], memory[29486], memory[29487]};
wire [31:0] memory29488 = {memory[29488], memory[29489], memory[29490], memory[29491]};
wire [31:0] memory29492 = {memory[29492], memory[29493], memory[29494], memory[29495]};
wire [31:0] memory29496 = {memory[29496], memory[29497], memory[29498], memory[29499]};
wire [31:0] memory29500 = {memory[29500], memory[29501], memory[29502], memory[29503]};
wire [31:0] memory29504 = {memory[29504], memory[29505], memory[29506], memory[29507]};
wire [31:0] memory29508 = {memory[29508], memory[29509], memory[29510], memory[29511]};
wire [31:0] memory29512 = {memory[29512], memory[29513], memory[29514], memory[29515]};
wire [31:0] memory29516 = {memory[29516], memory[29517], memory[29518], memory[29519]};
wire [31:0] memory29520 = {memory[29520], memory[29521], memory[29522], memory[29523]};
wire [31:0] memory29524 = {memory[29524], memory[29525], memory[29526], memory[29527]};
wire [31:0] memory29528 = {memory[29528], memory[29529], memory[29530], memory[29531]};
wire [31:0] memory29532 = {memory[29532], memory[29533], memory[29534], memory[29535]};
wire [31:0] memory29536 = {memory[29536], memory[29537], memory[29538], memory[29539]};
wire [31:0] memory29540 = {memory[29540], memory[29541], memory[29542], memory[29543]};
wire [31:0] memory29544 = {memory[29544], memory[29545], memory[29546], memory[29547]};
wire [31:0] memory29548 = {memory[29548], memory[29549], memory[29550], memory[29551]};
wire [31:0] memory29552 = {memory[29552], memory[29553], memory[29554], memory[29555]};
wire [31:0] memory29556 = {memory[29556], memory[29557], memory[29558], memory[29559]};
wire [31:0] memory29560 = {memory[29560], memory[29561], memory[29562], memory[29563]};
wire [31:0] memory29564 = {memory[29564], memory[29565], memory[29566], memory[29567]};
wire [31:0] memory29568 = {memory[29568], memory[29569], memory[29570], memory[29571]};
wire [31:0] memory29572 = {memory[29572], memory[29573], memory[29574], memory[29575]};
wire [31:0] memory29576 = {memory[29576], memory[29577], memory[29578], memory[29579]};
wire [31:0] memory29580 = {memory[29580], memory[29581], memory[29582], memory[29583]};
wire [31:0] memory29584 = {memory[29584], memory[29585], memory[29586], memory[29587]};
wire [31:0] memory29588 = {memory[29588], memory[29589], memory[29590], memory[29591]};
wire [31:0] memory29592 = {memory[29592], memory[29593], memory[29594], memory[29595]};
wire [31:0] memory29596 = {memory[29596], memory[29597], memory[29598], memory[29599]};
wire [31:0] memory29600 = {memory[29600], memory[29601], memory[29602], memory[29603]};
wire [31:0] memory29604 = {memory[29604], memory[29605], memory[29606], memory[29607]};
wire [31:0] memory29608 = {memory[29608], memory[29609], memory[29610], memory[29611]};
wire [31:0] memory29612 = {memory[29612], memory[29613], memory[29614], memory[29615]};
wire [31:0] memory29616 = {memory[29616], memory[29617], memory[29618], memory[29619]};
wire [31:0] memory29620 = {memory[29620], memory[29621], memory[29622], memory[29623]};
wire [31:0] memory29624 = {memory[29624], memory[29625], memory[29626], memory[29627]};
wire [31:0] memory29628 = {memory[29628], memory[29629], memory[29630], memory[29631]};
wire [31:0] memory29632 = {memory[29632], memory[29633], memory[29634], memory[29635]};
wire [31:0] memory29636 = {memory[29636], memory[29637], memory[29638], memory[29639]};
wire [31:0] memory29640 = {memory[29640], memory[29641], memory[29642], memory[29643]};
wire [31:0] memory29644 = {memory[29644], memory[29645], memory[29646], memory[29647]};
wire [31:0] memory29648 = {memory[29648], memory[29649], memory[29650], memory[29651]};
wire [31:0] memory29652 = {memory[29652], memory[29653], memory[29654], memory[29655]};
wire [31:0] memory29656 = {memory[29656], memory[29657], memory[29658], memory[29659]};
wire [31:0] memory29660 = {memory[29660], memory[29661], memory[29662], memory[29663]};
wire [31:0] memory29664 = {memory[29664], memory[29665], memory[29666], memory[29667]};
wire [31:0] memory29668 = {memory[29668], memory[29669], memory[29670], memory[29671]};
wire [31:0] memory29672 = {memory[29672], memory[29673], memory[29674], memory[29675]};
wire [31:0] memory29676 = {memory[29676], memory[29677], memory[29678], memory[29679]};
wire [31:0] memory29680 = {memory[29680], memory[29681], memory[29682], memory[29683]};
wire [31:0] memory29684 = {memory[29684], memory[29685], memory[29686], memory[29687]};
wire [31:0] memory29688 = {memory[29688], memory[29689], memory[29690], memory[29691]};
wire [31:0] memory29692 = {memory[29692], memory[29693], memory[29694], memory[29695]};
wire [31:0] memory29696 = {memory[29696], memory[29697], memory[29698], memory[29699]};
wire [31:0] memory29700 = {memory[29700], memory[29701], memory[29702], memory[29703]};
wire [31:0] memory29704 = {memory[29704], memory[29705], memory[29706], memory[29707]};
wire [31:0] memory29708 = {memory[29708], memory[29709], memory[29710], memory[29711]};
wire [31:0] memory29712 = {memory[29712], memory[29713], memory[29714], memory[29715]};
wire [31:0] memory29716 = {memory[29716], memory[29717], memory[29718], memory[29719]};
wire [31:0] memory29720 = {memory[29720], memory[29721], memory[29722], memory[29723]};
wire [31:0] memory29724 = {memory[29724], memory[29725], memory[29726], memory[29727]};
wire [31:0] memory29728 = {memory[29728], memory[29729], memory[29730], memory[29731]};
wire [31:0] memory29732 = {memory[29732], memory[29733], memory[29734], memory[29735]};
wire [31:0] memory29736 = {memory[29736], memory[29737], memory[29738], memory[29739]};
wire [31:0] memory29740 = {memory[29740], memory[29741], memory[29742], memory[29743]};
wire [31:0] memory29744 = {memory[29744], memory[29745], memory[29746], memory[29747]};
wire [31:0] memory29748 = {memory[29748], memory[29749], memory[29750], memory[29751]};
wire [31:0] memory29752 = {memory[29752], memory[29753], memory[29754], memory[29755]};
wire [31:0] memory29756 = {memory[29756], memory[29757], memory[29758], memory[29759]};
wire [31:0] memory29760 = {memory[29760], memory[29761], memory[29762], memory[29763]};
wire [31:0] memory29764 = {memory[29764], memory[29765], memory[29766], memory[29767]};
wire [31:0] memory29768 = {memory[29768], memory[29769], memory[29770], memory[29771]};
wire [31:0] memory29772 = {memory[29772], memory[29773], memory[29774], memory[29775]};
wire [31:0] memory29776 = {memory[29776], memory[29777], memory[29778], memory[29779]};
wire [31:0] memory29780 = {memory[29780], memory[29781], memory[29782], memory[29783]};
wire [31:0] memory29784 = {memory[29784], memory[29785], memory[29786], memory[29787]};
wire [31:0] memory29788 = {memory[29788], memory[29789], memory[29790], memory[29791]};
wire [31:0] memory29792 = {memory[29792], memory[29793], memory[29794], memory[29795]};
wire [31:0] memory29796 = {memory[29796], memory[29797], memory[29798], memory[29799]};
wire [31:0] memory29800 = {memory[29800], memory[29801], memory[29802], memory[29803]};
wire [31:0] memory29804 = {memory[29804], memory[29805], memory[29806], memory[29807]};
wire [31:0] memory29808 = {memory[29808], memory[29809], memory[29810], memory[29811]};
wire [31:0] memory29812 = {memory[29812], memory[29813], memory[29814], memory[29815]};
wire [31:0] memory29816 = {memory[29816], memory[29817], memory[29818], memory[29819]};
wire [31:0] memory29820 = {memory[29820], memory[29821], memory[29822], memory[29823]};
wire [31:0] memory29824 = {memory[29824], memory[29825], memory[29826], memory[29827]};
wire [31:0] memory29828 = {memory[29828], memory[29829], memory[29830], memory[29831]};
wire [31:0] memory29832 = {memory[29832], memory[29833], memory[29834], memory[29835]};
wire [31:0] memory29836 = {memory[29836], memory[29837], memory[29838], memory[29839]};
wire [31:0] memory29840 = {memory[29840], memory[29841], memory[29842], memory[29843]};
wire [31:0] memory29844 = {memory[29844], memory[29845], memory[29846], memory[29847]};
wire [31:0] memory29848 = {memory[29848], memory[29849], memory[29850], memory[29851]};
wire [31:0] memory29852 = {memory[29852], memory[29853], memory[29854], memory[29855]};
wire [31:0] memory29856 = {memory[29856], memory[29857], memory[29858], memory[29859]};
wire [31:0] memory29860 = {memory[29860], memory[29861], memory[29862], memory[29863]};
wire [31:0] memory29864 = {memory[29864], memory[29865], memory[29866], memory[29867]};
wire [31:0] memory29868 = {memory[29868], memory[29869], memory[29870], memory[29871]};
wire [31:0] memory29872 = {memory[29872], memory[29873], memory[29874], memory[29875]};
wire [31:0] memory29876 = {memory[29876], memory[29877], memory[29878], memory[29879]};
wire [31:0] memory29880 = {memory[29880], memory[29881], memory[29882], memory[29883]};
wire [31:0] memory29884 = {memory[29884], memory[29885], memory[29886], memory[29887]};
wire [31:0] memory29888 = {memory[29888], memory[29889], memory[29890], memory[29891]};
wire [31:0] memory29892 = {memory[29892], memory[29893], memory[29894], memory[29895]};
wire [31:0] memory29896 = {memory[29896], memory[29897], memory[29898], memory[29899]};
wire [31:0] memory29900 = {memory[29900], memory[29901], memory[29902], memory[29903]};
wire [31:0] memory29904 = {memory[29904], memory[29905], memory[29906], memory[29907]};
wire [31:0] memory29908 = {memory[29908], memory[29909], memory[29910], memory[29911]};
wire [31:0] memory29912 = {memory[29912], memory[29913], memory[29914], memory[29915]};
wire [31:0] memory29916 = {memory[29916], memory[29917], memory[29918], memory[29919]};
wire [31:0] memory29920 = {memory[29920], memory[29921], memory[29922], memory[29923]};
wire [31:0] memory29924 = {memory[29924], memory[29925], memory[29926], memory[29927]};
wire [31:0] memory29928 = {memory[29928], memory[29929], memory[29930], memory[29931]};
wire [31:0] memory29932 = {memory[29932], memory[29933], memory[29934], memory[29935]};
wire [31:0] memory29936 = {memory[29936], memory[29937], memory[29938], memory[29939]};
wire [31:0] memory29940 = {memory[29940], memory[29941], memory[29942], memory[29943]};
wire [31:0] memory29944 = {memory[29944], memory[29945], memory[29946], memory[29947]};
wire [31:0] memory29948 = {memory[29948], memory[29949], memory[29950], memory[29951]};
wire [31:0] memory29952 = {memory[29952], memory[29953], memory[29954], memory[29955]};
wire [31:0] memory29956 = {memory[29956], memory[29957], memory[29958], memory[29959]};
wire [31:0] memory29960 = {memory[29960], memory[29961], memory[29962], memory[29963]};
wire [31:0] memory29964 = {memory[29964], memory[29965], memory[29966], memory[29967]};
wire [31:0] memory29968 = {memory[29968], memory[29969], memory[29970], memory[29971]};
wire [31:0] memory29972 = {memory[29972], memory[29973], memory[29974], memory[29975]};
wire [31:0] memory29976 = {memory[29976], memory[29977], memory[29978], memory[29979]};
wire [31:0] memory29980 = {memory[29980], memory[29981], memory[29982], memory[29983]};
wire [31:0] memory29984 = {memory[29984], memory[29985], memory[29986], memory[29987]};
wire [31:0] memory29988 = {memory[29988], memory[29989], memory[29990], memory[29991]};
wire [31:0] memory29992 = {memory[29992], memory[29993], memory[29994], memory[29995]};
wire [31:0] memory29996 = {memory[29996], memory[29997], memory[29998], memory[29999]};
wire [31:0] memory30000 = {memory[30000], memory[30001], memory[30002], memory[30003]};
wire [31:0] memory30004 = {memory[30004], memory[30005], memory[30006], memory[30007]};
wire [31:0] memory30008 = {memory[30008], memory[30009], memory[30010], memory[30011]};
wire [31:0] memory30012 = {memory[30012], memory[30013], memory[30014], memory[30015]};
wire [31:0] memory30016 = {memory[30016], memory[30017], memory[30018], memory[30019]};
wire [31:0] memory30020 = {memory[30020], memory[30021], memory[30022], memory[30023]};
wire [31:0] memory30024 = {memory[30024], memory[30025], memory[30026], memory[30027]};
wire [31:0] memory30028 = {memory[30028], memory[30029], memory[30030], memory[30031]};
wire [31:0] memory30032 = {memory[30032], memory[30033], memory[30034], memory[30035]};
wire [31:0] memory30036 = {memory[30036], memory[30037], memory[30038], memory[30039]};
wire [31:0] memory30040 = {memory[30040], memory[30041], memory[30042], memory[30043]};
wire [31:0] memory30044 = {memory[30044], memory[30045], memory[30046], memory[30047]};
wire [31:0] memory30048 = {memory[30048], memory[30049], memory[30050], memory[30051]};
wire [31:0] memory30052 = {memory[30052], memory[30053], memory[30054], memory[30055]};
wire [31:0] memory30056 = {memory[30056], memory[30057], memory[30058], memory[30059]};
wire [31:0] memory30060 = {memory[30060], memory[30061], memory[30062], memory[30063]};
wire [31:0] memory30064 = {memory[30064], memory[30065], memory[30066], memory[30067]};
wire [31:0] memory30068 = {memory[30068], memory[30069], memory[30070], memory[30071]};
wire [31:0] memory30072 = {memory[30072], memory[30073], memory[30074], memory[30075]};
wire [31:0] memory30076 = {memory[30076], memory[30077], memory[30078], memory[30079]};
wire [31:0] memory30080 = {memory[30080], memory[30081], memory[30082], memory[30083]};
wire [31:0] memory30084 = {memory[30084], memory[30085], memory[30086], memory[30087]};
wire [31:0] memory30088 = {memory[30088], memory[30089], memory[30090], memory[30091]};
wire [31:0] memory30092 = {memory[30092], memory[30093], memory[30094], memory[30095]};
wire [31:0] memory30096 = {memory[30096], memory[30097], memory[30098], memory[30099]};
wire [31:0] memory30100 = {memory[30100], memory[30101], memory[30102], memory[30103]};
wire [31:0] memory30104 = {memory[30104], memory[30105], memory[30106], memory[30107]};
wire [31:0] memory30108 = {memory[30108], memory[30109], memory[30110], memory[30111]};
wire [31:0] memory30112 = {memory[30112], memory[30113], memory[30114], memory[30115]};
wire [31:0] memory30116 = {memory[30116], memory[30117], memory[30118], memory[30119]};
wire [31:0] memory30120 = {memory[30120], memory[30121], memory[30122], memory[30123]};
wire [31:0] memory30124 = {memory[30124], memory[30125], memory[30126], memory[30127]};
wire [31:0] memory30128 = {memory[30128], memory[30129], memory[30130], memory[30131]};
wire [31:0] memory30132 = {memory[30132], memory[30133], memory[30134], memory[30135]};
wire [31:0] memory30136 = {memory[30136], memory[30137], memory[30138], memory[30139]};
wire [31:0] memory30140 = {memory[30140], memory[30141], memory[30142], memory[30143]};
wire [31:0] memory30144 = {memory[30144], memory[30145], memory[30146], memory[30147]};
wire [31:0] memory30148 = {memory[30148], memory[30149], memory[30150], memory[30151]};
wire [31:0] memory30152 = {memory[30152], memory[30153], memory[30154], memory[30155]};
wire [31:0] memory30156 = {memory[30156], memory[30157], memory[30158], memory[30159]};
wire [31:0] memory30160 = {memory[30160], memory[30161], memory[30162], memory[30163]};
wire [31:0] memory30164 = {memory[30164], memory[30165], memory[30166], memory[30167]};
wire [31:0] memory30168 = {memory[30168], memory[30169], memory[30170], memory[30171]};
wire [31:0] memory30172 = {memory[30172], memory[30173], memory[30174], memory[30175]};
wire [31:0] memory30176 = {memory[30176], memory[30177], memory[30178], memory[30179]};
wire [31:0] memory30180 = {memory[30180], memory[30181], memory[30182], memory[30183]};
wire [31:0] memory30184 = {memory[30184], memory[30185], memory[30186], memory[30187]};
wire [31:0] memory30188 = {memory[30188], memory[30189], memory[30190], memory[30191]};
wire [31:0] memory30192 = {memory[30192], memory[30193], memory[30194], memory[30195]};
wire [31:0] memory30196 = {memory[30196], memory[30197], memory[30198], memory[30199]};
wire [31:0] memory30200 = {memory[30200], memory[30201], memory[30202], memory[30203]};
wire [31:0] memory30204 = {memory[30204], memory[30205], memory[30206], memory[30207]};
wire [31:0] memory30208 = {memory[30208], memory[30209], memory[30210], memory[30211]};
wire [31:0] memory30212 = {memory[30212], memory[30213], memory[30214], memory[30215]};
wire [31:0] memory30216 = {memory[30216], memory[30217], memory[30218], memory[30219]};
wire [31:0] memory30220 = {memory[30220], memory[30221], memory[30222], memory[30223]};
wire [31:0] memory30224 = {memory[30224], memory[30225], memory[30226], memory[30227]};
wire [31:0] memory30228 = {memory[30228], memory[30229], memory[30230], memory[30231]};
wire [31:0] memory30232 = {memory[30232], memory[30233], memory[30234], memory[30235]};
wire [31:0] memory30236 = {memory[30236], memory[30237], memory[30238], memory[30239]};
wire [31:0] memory30240 = {memory[30240], memory[30241], memory[30242], memory[30243]};
wire [31:0] memory30244 = {memory[30244], memory[30245], memory[30246], memory[30247]};
wire [31:0] memory30248 = {memory[30248], memory[30249], memory[30250], memory[30251]};
wire [31:0] memory30252 = {memory[30252], memory[30253], memory[30254], memory[30255]};
wire [31:0] memory30256 = {memory[30256], memory[30257], memory[30258], memory[30259]};
wire [31:0] memory30260 = {memory[30260], memory[30261], memory[30262], memory[30263]};
wire [31:0] memory30264 = {memory[30264], memory[30265], memory[30266], memory[30267]};
wire [31:0] memory30268 = {memory[30268], memory[30269], memory[30270], memory[30271]};
wire [31:0] memory30272 = {memory[30272], memory[30273], memory[30274], memory[30275]};
wire [31:0] memory30276 = {memory[30276], memory[30277], memory[30278], memory[30279]};
wire [31:0] memory30280 = {memory[30280], memory[30281], memory[30282], memory[30283]};
wire [31:0] memory30284 = {memory[30284], memory[30285], memory[30286], memory[30287]};
wire [31:0] memory30288 = {memory[30288], memory[30289], memory[30290], memory[30291]};
wire [31:0] memory30292 = {memory[30292], memory[30293], memory[30294], memory[30295]};
wire [31:0] memory30296 = {memory[30296], memory[30297], memory[30298], memory[30299]};
wire [31:0] memory30300 = {memory[30300], memory[30301], memory[30302], memory[30303]};
wire [31:0] memory30304 = {memory[30304], memory[30305], memory[30306], memory[30307]};
wire [31:0] memory30308 = {memory[30308], memory[30309], memory[30310], memory[30311]};
wire [31:0] memory30312 = {memory[30312], memory[30313], memory[30314], memory[30315]};
wire [31:0] memory30316 = {memory[30316], memory[30317], memory[30318], memory[30319]};
wire [31:0] memory30320 = {memory[30320], memory[30321], memory[30322], memory[30323]};
wire [31:0] memory30324 = {memory[30324], memory[30325], memory[30326], memory[30327]};
wire [31:0] memory30328 = {memory[30328], memory[30329], memory[30330], memory[30331]};
wire [31:0] memory30332 = {memory[30332], memory[30333], memory[30334], memory[30335]};
wire [31:0] memory30336 = {memory[30336], memory[30337], memory[30338], memory[30339]};
wire [31:0] memory30340 = {memory[30340], memory[30341], memory[30342], memory[30343]};
wire [31:0] memory30344 = {memory[30344], memory[30345], memory[30346], memory[30347]};
wire [31:0] memory30348 = {memory[30348], memory[30349], memory[30350], memory[30351]};
wire [31:0] memory30352 = {memory[30352], memory[30353], memory[30354], memory[30355]};
wire [31:0] memory30356 = {memory[30356], memory[30357], memory[30358], memory[30359]};
wire [31:0] memory30360 = {memory[30360], memory[30361], memory[30362], memory[30363]};
wire [31:0] memory30364 = {memory[30364], memory[30365], memory[30366], memory[30367]};
wire [31:0] memory30368 = {memory[30368], memory[30369], memory[30370], memory[30371]};
wire [31:0] memory30372 = {memory[30372], memory[30373], memory[30374], memory[30375]};
wire [31:0] memory30376 = {memory[30376], memory[30377], memory[30378], memory[30379]};
wire [31:0] memory30380 = {memory[30380], memory[30381], memory[30382], memory[30383]};
wire [31:0] memory30384 = {memory[30384], memory[30385], memory[30386], memory[30387]};
wire [31:0] memory30388 = {memory[30388], memory[30389], memory[30390], memory[30391]};
wire [31:0] memory30392 = {memory[30392], memory[30393], memory[30394], memory[30395]};
wire [31:0] memory30396 = {memory[30396], memory[30397], memory[30398], memory[30399]};
wire [31:0] memory30400 = {memory[30400], memory[30401], memory[30402], memory[30403]};
wire [31:0] memory30404 = {memory[30404], memory[30405], memory[30406], memory[30407]};
wire [31:0] memory30408 = {memory[30408], memory[30409], memory[30410], memory[30411]};
wire [31:0] memory30412 = {memory[30412], memory[30413], memory[30414], memory[30415]};
wire [31:0] memory30416 = {memory[30416], memory[30417], memory[30418], memory[30419]};
wire [31:0] memory30420 = {memory[30420], memory[30421], memory[30422], memory[30423]};
wire [31:0] memory30424 = {memory[30424], memory[30425], memory[30426], memory[30427]};
wire [31:0] memory30428 = {memory[30428], memory[30429], memory[30430], memory[30431]};
wire [31:0] memory30432 = {memory[30432], memory[30433], memory[30434], memory[30435]};
wire [31:0] memory30436 = {memory[30436], memory[30437], memory[30438], memory[30439]};
wire [31:0] memory30440 = {memory[30440], memory[30441], memory[30442], memory[30443]};
wire [31:0] memory30444 = {memory[30444], memory[30445], memory[30446], memory[30447]};
wire [31:0] memory30448 = {memory[30448], memory[30449], memory[30450], memory[30451]};
wire [31:0] memory30452 = {memory[30452], memory[30453], memory[30454], memory[30455]};
wire [31:0] memory30456 = {memory[30456], memory[30457], memory[30458], memory[30459]};
wire [31:0] memory30460 = {memory[30460], memory[30461], memory[30462], memory[30463]};
wire [31:0] memory30464 = {memory[30464], memory[30465], memory[30466], memory[30467]};
wire [31:0] memory30468 = {memory[30468], memory[30469], memory[30470], memory[30471]};
wire [31:0] memory30472 = {memory[30472], memory[30473], memory[30474], memory[30475]};
wire [31:0] memory30476 = {memory[30476], memory[30477], memory[30478], memory[30479]};
wire [31:0] memory30480 = {memory[30480], memory[30481], memory[30482], memory[30483]};
wire [31:0] memory30484 = {memory[30484], memory[30485], memory[30486], memory[30487]};
wire [31:0] memory30488 = {memory[30488], memory[30489], memory[30490], memory[30491]};
wire [31:0] memory30492 = {memory[30492], memory[30493], memory[30494], memory[30495]};
wire [31:0] memory30496 = {memory[30496], memory[30497], memory[30498], memory[30499]};
wire [31:0] memory30500 = {memory[30500], memory[30501], memory[30502], memory[30503]};
wire [31:0] memory30504 = {memory[30504], memory[30505], memory[30506], memory[30507]};
wire [31:0] memory30508 = {memory[30508], memory[30509], memory[30510], memory[30511]};
wire [31:0] memory30512 = {memory[30512], memory[30513], memory[30514], memory[30515]};
wire [31:0] memory30516 = {memory[30516], memory[30517], memory[30518], memory[30519]};
wire [31:0] memory30520 = {memory[30520], memory[30521], memory[30522], memory[30523]};
wire [31:0] memory30524 = {memory[30524], memory[30525], memory[30526], memory[30527]};
wire [31:0] memory30528 = {memory[30528], memory[30529], memory[30530], memory[30531]};
wire [31:0] memory30532 = {memory[30532], memory[30533], memory[30534], memory[30535]};
wire [31:0] memory30536 = {memory[30536], memory[30537], memory[30538], memory[30539]};
wire [31:0] memory30540 = {memory[30540], memory[30541], memory[30542], memory[30543]};
wire [31:0] memory30544 = {memory[30544], memory[30545], memory[30546], memory[30547]};
wire [31:0] memory30548 = {memory[30548], memory[30549], memory[30550], memory[30551]};
wire [31:0] memory30552 = {memory[30552], memory[30553], memory[30554], memory[30555]};
wire [31:0] memory30556 = {memory[30556], memory[30557], memory[30558], memory[30559]};
wire [31:0] memory30560 = {memory[30560], memory[30561], memory[30562], memory[30563]};
wire [31:0] memory30564 = {memory[30564], memory[30565], memory[30566], memory[30567]};
wire [31:0] memory30568 = {memory[30568], memory[30569], memory[30570], memory[30571]};
wire [31:0] memory30572 = {memory[30572], memory[30573], memory[30574], memory[30575]};
wire [31:0] memory30576 = {memory[30576], memory[30577], memory[30578], memory[30579]};
wire [31:0] memory30580 = {memory[30580], memory[30581], memory[30582], memory[30583]};
wire [31:0] memory30584 = {memory[30584], memory[30585], memory[30586], memory[30587]};
wire [31:0] memory30588 = {memory[30588], memory[30589], memory[30590], memory[30591]};
wire [31:0] memory30592 = {memory[30592], memory[30593], memory[30594], memory[30595]};
wire [31:0] memory30596 = {memory[30596], memory[30597], memory[30598], memory[30599]};
wire [31:0] memory30600 = {memory[30600], memory[30601], memory[30602], memory[30603]};
wire [31:0] memory30604 = {memory[30604], memory[30605], memory[30606], memory[30607]};
wire [31:0] memory30608 = {memory[30608], memory[30609], memory[30610], memory[30611]};
wire [31:0] memory30612 = {memory[30612], memory[30613], memory[30614], memory[30615]};
wire [31:0] memory30616 = {memory[30616], memory[30617], memory[30618], memory[30619]};
wire [31:0] memory30620 = {memory[30620], memory[30621], memory[30622], memory[30623]};
wire [31:0] memory30624 = {memory[30624], memory[30625], memory[30626], memory[30627]};
wire [31:0] memory30628 = {memory[30628], memory[30629], memory[30630], memory[30631]};
wire [31:0] memory30632 = {memory[30632], memory[30633], memory[30634], memory[30635]};
wire [31:0] memory30636 = {memory[30636], memory[30637], memory[30638], memory[30639]};
wire [31:0] memory30640 = {memory[30640], memory[30641], memory[30642], memory[30643]};
wire [31:0] memory30644 = {memory[30644], memory[30645], memory[30646], memory[30647]};
wire [31:0] memory30648 = {memory[30648], memory[30649], memory[30650], memory[30651]};
wire [31:0] memory30652 = {memory[30652], memory[30653], memory[30654], memory[30655]};
wire [31:0] memory30656 = {memory[30656], memory[30657], memory[30658], memory[30659]};
wire [31:0] memory30660 = {memory[30660], memory[30661], memory[30662], memory[30663]};
wire [31:0] memory30664 = {memory[30664], memory[30665], memory[30666], memory[30667]};
wire [31:0] memory30668 = {memory[30668], memory[30669], memory[30670], memory[30671]};
wire [31:0] memory30672 = {memory[30672], memory[30673], memory[30674], memory[30675]};
wire [31:0] memory30676 = {memory[30676], memory[30677], memory[30678], memory[30679]};
wire [31:0] memory30680 = {memory[30680], memory[30681], memory[30682], memory[30683]};
wire [31:0] memory30684 = {memory[30684], memory[30685], memory[30686], memory[30687]};
wire [31:0] memory30688 = {memory[30688], memory[30689], memory[30690], memory[30691]};
wire [31:0] memory30692 = {memory[30692], memory[30693], memory[30694], memory[30695]};
wire [31:0] memory30696 = {memory[30696], memory[30697], memory[30698], memory[30699]};
wire [31:0] memory30700 = {memory[30700], memory[30701], memory[30702], memory[30703]};
wire [31:0] memory30704 = {memory[30704], memory[30705], memory[30706], memory[30707]};
wire [31:0] memory30708 = {memory[30708], memory[30709], memory[30710], memory[30711]};
wire [31:0] memory30712 = {memory[30712], memory[30713], memory[30714], memory[30715]};

endmodule
